magic
tech sky130A
magscale 1 2
timestamp 1739975917
<< locali >>
rect 1013 468 2229 506
rect 1013 413 1667 468
rect 1013 -720 1098 413
rect 1546 316 1667 413
rect 1992 316 2229 468
rect 1546 4 2229 316
rect 1546 -100 1697 4
rect 1751 -100 2229 4
rect 1546 -189 2229 -100
rect 1546 -720 1690 -189
rect 2138 -720 2229 -189
rect 1012 -2164 1097 -1050
rect 1545 -1564 1689 -1050
rect 2135 -1564 2229 -1050
rect 1545 -1620 2229 -1564
rect 1545 -1729 1696 -1620
rect 1755 -1729 2229 -1620
rect 1545 -2062 2229 -1729
rect 1545 -2164 1667 -2062
rect 1012 -2230 1667 -2164
rect 1990 -2230 2229 -2062
rect 1012 -2269 2229 -2230
<< viali >>
rect 1667 316 1992 468
rect 1697 -100 1751 4
rect 1696 -1729 1755 -1620
rect 1667 -2230 1990 -2062
<< metal1 >>
rect 1638 468 2214 489
rect 1149 -521 1159 -136
rect 1211 -521 1221 -136
rect 1291 -796 1351 347
rect 1638 316 1667 468
rect 1992 316 2214 468
rect 1638 289 2214 316
rect 1678 -109 1688 11
rect 1759 -109 1769 11
rect 1424 -523 1434 -139
rect 1494 -523 1504 -139
rect 1738 -520 1748 -349
rect 1800 -520 1810 -349
rect 1290 -862 1351 -796
rect 1883 -847 1943 -253
rect 2017 -521 2027 -349
rect 2081 -521 2091 -349
rect 1732 -852 1943 -847
rect 1272 -866 1351 -862
rect 1268 -918 1278 -866
rect 1340 -918 1351 -866
rect 1272 -922 1351 -918
rect 1728 -921 1738 -852
rect 1794 -921 1943 -852
rect 1290 -988 1351 -922
rect 1732 -927 1943 -921
rect 1149 -1616 1159 -1237
rect 1211 -1616 1221 -1237
rect 1291 -2099 1351 -988
rect 1425 -1622 1435 -1238
rect 1495 -1622 1505 -1238
rect 1737 -1412 1747 -1240
rect 1799 -1412 1809 -1240
rect 1883 -1499 1943 -927
rect 2018 -1408 2028 -1242
rect 2082 -1408 2092 -1242
rect 1679 -1735 1689 -1612
rect 1761 -1735 1771 -1612
rect 1647 -2062 2208 -2047
rect 1647 -2230 1667 -2062
rect 1990 -2230 2208 -2062
rect 1647 -2247 2208 -2230
<< via1 >>
rect 1159 -521 1211 -136
rect 1688 4 1759 11
rect 1688 -100 1697 4
rect 1697 -100 1751 4
rect 1751 -100 1759 4
rect 1688 -109 1759 -100
rect 1434 -523 1494 -139
rect 1748 -520 1800 -349
rect 2027 -521 2081 -349
rect 1278 -918 1340 -866
rect 1738 -921 1794 -852
rect 1159 -1616 1211 -1237
rect 1435 -1622 1495 -1238
rect 1747 -1412 1799 -1240
rect 2028 -1408 2082 -1242
rect 1689 -1620 1761 -1612
rect 1689 -1729 1696 -1620
rect 1696 -1729 1755 -1620
rect 1755 -1729 1761 -1620
rect 1689 -1735 1761 -1729
<< metal2 >>
rect 1688 16 1759 21
rect 1682 11 1765 16
rect 1682 -109 1688 11
rect 1759 -109 1765 11
rect 1159 -133 1211 -126
rect 1149 -136 1211 -133
rect 1149 -393 1159 -136
rect 1013 -521 1159 -393
rect 1434 -137 1494 -129
rect 1432 -139 1551 -137
rect 1211 -521 1215 -393
rect 1013 -593 1215 -521
rect 1432 -523 1434 -139
rect 1494 -523 1551 -139
rect 1432 -525 1551 -523
rect 1682 -339 1765 -109
rect 1682 -346 1800 -339
rect 2027 -346 2081 -339
rect 1682 -349 1803 -346
rect 1682 -520 1748 -349
rect 1800 -520 1803 -349
rect 1682 -524 1803 -520
rect 2024 -349 2146 -346
rect 2024 -521 2027 -349
rect 2081 -521 2146 -349
rect 2024 -524 2146 -521
rect 1434 -533 1551 -525
rect 1748 -530 1800 -524
rect 2027 -531 2146 -524
rect 1146 -866 1346 -792
rect 1146 -918 1278 -866
rect 1340 -918 1346 -866
rect 1146 -992 1346 -918
rect 1480 -847 1551 -533
rect 2065 -792 2146 -531
rect 1738 -847 1794 -842
rect 1480 -852 1799 -847
rect 1480 -921 1738 -852
rect 1794 -921 1799 -852
rect 1480 -927 1799 -921
rect 1012 -1237 1214 -1166
rect 1480 -1228 1551 -927
rect 1738 -931 1794 -927
rect 2064 -992 2266 -792
rect 1435 -1236 1551 -1228
rect 1012 -1366 1159 -1237
rect 1149 -1616 1159 -1366
rect 1211 -1366 1214 -1237
rect 1432 -1238 1551 -1236
rect 1747 -1237 1799 -1230
rect 2065 -1232 2146 -992
rect 2028 -1236 2146 -1232
rect 1149 -1623 1211 -1616
rect 1159 -1626 1211 -1623
rect 1432 -1622 1435 -1238
rect 1495 -1622 1551 -1238
rect 1432 -1625 1551 -1622
rect 1683 -1240 1802 -1237
rect 1683 -1412 1747 -1240
rect 1799 -1412 1802 -1240
rect 1683 -1415 1802 -1412
rect 2024 -1242 2146 -1236
rect 2024 -1408 2028 -1242
rect 2082 -1408 2146 -1242
rect 2024 -1415 2146 -1408
rect 1683 -1422 1799 -1415
rect 2028 -1418 2082 -1415
rect 1683 -1612 1766 -1422
rect 1435 -1632 1495 -1625
rect 1683 -1735 1689 -1612
rect 1761 -1735 1766 -1612
rect 1683 -1741 1766 -1735
rect 1689 -1745 1761 -1741
use sky130_fd_pr__pfet_01v8_lvt_3VA8VM  XM1
timestamp 1739902357
transform 1 0 1322 0 1 -134
box -296 -619 296 619
use sky130_fd_pr__nfet_01v8_lvt_AHMAL2  XM2
timestamp 1739797948
transform -1 0 1321 0 1 -1625
box -296 -610 296 610
use sky130_fd_pr__pfet_01v8_lvt_3VR9VM  XM3
timestamp 1739797948
transform 1 0 1914 0 1 -434
box -296 -319 296 319
use sky130_fd_pr__nfet_01v8_lvt_69TQ3K  XM4
timestamp 1739797948
transform 1 0 1913 0 1 -1325
box -296 -310 296 310
<< labels >>
flabel metal1 2014 289 2214 489 0 FreeSans 256 0 0 0 VPWR
port 0 nsew
flabel metal1 2008 -2247 2208 -2047 0 FreeSans 256 0 0 0 VGND
port 5 nsew
flabel metal2 2064 -992 2264 -792 0 FreeSans 256 0 0 0 Vcomp
port 3 nsew
flabel metal2 1146 -992 1346 -792 0 FreeSans 256 0 0 0 D3
port 2 nsew
flabel metal2 1012 -1366 1212 -1166 0 FreeSans 256 0 0 0 Vcomp_n
port 4 nsew
flabel metal2 1013 -593 1213 -393 0 FreeSans 256 0 0 0 Vcomp_p
port 1 nsew
<< end >>
