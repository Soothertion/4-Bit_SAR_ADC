magic
tech sky130A
timestamp 1740063090
<< poly >>
rect -700 500 -600 600
rect -100 500 400 600
rect 600 500 900 600
rect 1100 500 1600 600
rect 2200 500 2600 600
rect 3000 500 3100 600
rect 3400 500 3900 600
rect 4600 500 4700 600
rect 5000 500 5400 600
rect 5800 500 6100 600
rect -800 400 -600 500
rect -900 385 -785 400
rect -900 300 -800 385
rect -1000 285 -885 300
rect -1000 200 -900 285
rect -700 200 -600 400
rect 0 300 100 500
rect 385 485 500 500
rect 400 315 500 485
rect 385 300 500 315
rect -400 200 -200 300
rect 0 200 400 300
rect -1000 100 -500 200
rect -700 -100 -600 100
rect 0 0 100 200
rect 385 185 500 200
rect 400 15 500 185
rect 385 0 500 15
rect 700 0 800 500
rect 1000 485 1115 500
rect 1000 400 1100 485
rect 1300 0 1400 500
rect 1585 485 1700 500
rect 1600 400 1700 485
rect 2100 485 2215 500
rect 2585 485 2700 500
rect 2100 315 2200 485
rect 2600 400 2700 485
rect 2900 485 3015 500
rect 3085 485 3200 500
rect 2900 400 3000 485
rect 3100 400 3200 485
rect 2800 385 2915 400
rect 3185 385 3300 400
rect 2100 300 2215 315
rect 2200 200 2600 300
rect 2800 200 2900 385
rect 3200 200 3300 385
rect 2585 185 2700 200
rect 2100 15 2200 100
rect 2600 15 2700 185
rect 2100 0 2215 15
rect 2585 0 2700 15
rect 2800 100 3300 200
rect -100 -100 400 0
rect 600 -100 900 0
rect 1200 -100 1500 0
rect 2200 -100 2600 0
rect 2800 -100 2900 100
rect 3200 -100 3300 100
rect 3500 300 3600 500
rect 3885 485 4000 500
rect 3900 315 4000 485
rect 4500 485 4615 500
rect 4685 485 4800 500
rect 4500 400 4600 485
rect 4700 400 4800 485
rect 3885 300 4000 315
rect 4400 385 4515 400
rect 4785 385 4900 400
rect 3500 200 3900 300
rect 4400 200 4500 385
rect 4800 200 4900 385
rect 3500 0 3600 200
rect 3700 100 3800 200
rect 4400 100 4900 200
rect 3785 85 3900 100
rect 3800 0 3900 85
rect 3400 -100 3700 0
rect 3885 -15 4000 0
rect 3900 -100 4000 -15
rect 4400 -100 4500 100
rect 4800 -100 4900 100
rect 5100 0 5200 500
rect 5385 485 5500 500
rect 5400 400 5500 485
rect 5700 485 5815 500
rect 6085 485 6200 500
rect 5485 385 5600 400
rect 5500 15 5600 385
rect 5485 0 5600 15
rect 5700 15 5800 485
rect 6100 400 6200 485
rect 6100 15 6200 100
rect 5700 0 5815 15
rect 6085 0 6200 15
rect 5000 -100 5500 0
rect 5800 -100 6100 0
rect -1000 -300 -750 -250
rect -950 -400 -900 -300
rect -765 -315 -700 -300
rect -750 -385 -700 -315
rect -765 -400 -700 -385
rect -950 -450 -750 -400
rect -950 -550 -900 -450
rect -850 -500 -800 -450
rect -815 -515 -750 -500
rect -800 -550 -750 -515
rect -650 -535 -600 -250
rect -450 -500 -400 -250
rect -300 -300 -250 -250
rect -50 -300 50 -250
rect 100 -300 150 -250
rect 350 -300 450 -250
rect 500 -300 650 -250
rect 700 -300 750 -250
rect 950 -300 1050 -250
rect 1150 -300 1300 -250
rect 1600 -300 1750 -250
rect 1850 -300 1900 -250
rect 2100 -300 2200 -250
rect 2350 -300 2500 -250
rect 2550 -300 2700 -250
rect 2800 -300 2950 -250
rect 3050 -300 3300 -250
rect 3450 -300 3650 -250
rect 3750 -300 3950 -250
rect 4300 -285 4350 -250
rect 4299 -300 4351 -285
rect 4500 -300 4550 -250
rect 4750 -300 4850 -250
rect 4900 -300 5100 -250
rect 5400 -300 5600 -250
rect 5750 -300 6000 -250
rect 6150 -300 6350 -250
rect 6500 -285 6550 -250
rect 6499 -300 6551 -285
rect 6700 -300 6800 -250
rect 7000 -300 7100 -250
rect 7200 -300 7400 -250
rect -265 -315 -200 -300
rect -500 -535 -400 -500
rect -650 -550 -585 -535
rect -515 -550 -400 -535
rect -250 -350 -200 -315
rect -250 -400 -150 -350
rect -250 -550 -200 -400
rect -165 -415 -100 -400
rect -150 -450 -100 -415
rect -50 -450 0 -300
rect 135 -315 200 -300
rect -115 -465 0 -450
rect -100 -500 0 -465
rect -1000 -600 -850 -550
rect -765 -565 -700 -550
rect -750 -600 -700 -565
rect -600 -600 -500 -550
rect -450 -600 -350 -550
rect -300 -600 -150 -550
rect -50 -600 0 -500
rect 150 -350 200 -315
rect 150 -400 250 -350
rect 150 -550 200 -400
rect 235 -415 300 -400
rect 250 -450 300 -415
rect 350 -450 400 -300
rect 285 -465 400 -450
rect 300 -500 400 -465
rect 100 -600 250 -550
rect 350 -600 400 -500
rect 550 -550 600 -300
rect 735 -315 800 -300
rect 750 -350 800 -315
rect 750 -400 850 -350
rect 750 -550 800 -400
rect 835 -415 900 -400
rect 850 -450 900 -415
rect 950 -450 1000 -300
rect 885 -465 1000 -450
rect 900 -500 1000 -465
rect 500 -600 650 -550
rect 700 -600 850 -550
rect 950 -600 1000 -500
rect 1100 -315 1165 -300
rect 1285 -315 1350 -300
rect 1100 -535 1150 -315
rect 1300 -350 1350 -315
rect 1550 -315 1615 -300
rect 1735 -315 1800 -300
rect 1885 -315 1950 -300
rect 1250 -500 1350 -450
rect 1300 -535 1350 -500
rect 1100 -550 1165 -535
rect 1285 -550 1350 -535
rect 1550 -535 1600 -315
rect 1750 -535 1800 -315
rect 1550 -550 1615 -535
rect 1735 -550 1800 -535
rect 1900 -350 1950 -315
rect 1900 -400 2000 -350
rect 1900 -550 1950 -400
rect 1985 -415 2050 -400
rect 2000 -450 2050 -415
rect 2100 -450 2150 -300
rect 2035 -465 2150 -450
rect 2050 -500 2150 -465
rect 1150 -600 1300 -550
rect 1600 -600 1750 -550
rect 1850 -600 2000 -550
rect 2100 -600 2150 -500
rect 2400 -400 2450 -300
rect 2600 -400 2650 -300
rect 2400 -450 2650 -400
rect 2400 -550 2450 -450
rect 2600 -550 2650 -450
rect 2750 -315 2815 -300
rect 2935 -315 3000 -300
rect 2750 -535 2800 -315
rect 2950 -535 3000 -315
rect 2750 -550 2815 -535
rect 2935 -550 3000 -535
rect 3100 -400 3150 -300
rect 3285 -315 3350 -300
rect 3300 -385 3350 -315
rect 3285 -400 3350 -385
rect 3400 -315 3465 -300
rect 3700 -315 3765 -300
rect 3935 -315 4000 -300
rect 3400 -400 3450 -315
rect 3700 -385 3750 -315
rect 3950 -350 4000 -315
rect 4250 -315 4314 -300
rect 4336 -315 4400 -300
rect 4535 -315 4600 -300
rect 4250 -350 4300 -315
rect 4350 -350 4400 -315
rect 4550 -350 4600 -315
rect 4200 -365 4265 -350
rect 4385 -365 4450 -350
rect 3700 -400 3765 -385
rect 3100 -450 3300 -400
rect 3400 -450 3600 -400
rect 3750 -450 3950 -400
rect 4200 -450 4250 -365
rect 4400 -450 4450 -365
rect 3100 -550 3150 -450
rect 3400 -535 3450 -450
rect 3935 -465 4000 -450
rect 3700 -535 3750 -500
rect 3950 -535 4000 -465
rect 3400 -550 3465 -535
rect 3700 -550 3765 -535
rect 3935 -550 4000 -535
rect 4200 -500 4450 -450
rect 2350 -600 2500 -550
rect 2550 -600 2700 -550
rect 2800 -600 2950 -550
rect 3050 -600 3200 -550
rect 3450 -600 3650 -550
rect 3750 -600 3950 -550
rect 4200 -600 4250 -500
rect 4400 -600 4450 -500
rect 4550 -400 4650 -350
rect 4550 -550 4600 -400
rect 4635 -415 4700 -400
rect 4650 -450 4700 -415
rect 4750 -450 4800 -300
rect 4685 -465 4800 -450
rect 4700 -500 4800 -465
rect 4500 -600 4650 -550
rect 4750 -600 4800 -500
rect 4950 -550 5000 -300
rect 5085 -315 5150 -300
rect 5100 -350 5150 -315
rect 5135 -365 5200 -350
rect 5150 -535 5200 -365
rect 5135 -550 5200 -535
rect 5450 -550 5500 -300
rect 5585 -315 5650 -300
rect 5600 -350 5650 -315
rect 5635 -365 5700 -350
rect 5650 -535 5700 -365
rect 5635 -550 5700 -535
rect 5800 -400 5850 -300
rect 5985 -315 6050 -300
rect 6000 -385 6050 -315
rect 5985 -400 6050 -385
rect 6100 -315 6165 -300
rect 6450 -315 6514 -300
rect 6536 -315 6600 -300
rect 6100 -400 6150 -315
rect 6450 -350 6500 -315
rect 6550 -350 6600 -315
rect 6750 -350 6850 -300
rect 6950 -350 7050 -300
rect 6400 -365 6465 -350
rect 6585 -365 6650 -350
rect 5800 -450 6000 -400
rect 6100 -450 6300 -400
rect 6400 -450 6450 -365
rect 6600 -450 6650 -365
rect 5800 -550 5850 -450
rect 5900 -500 5950 -450
rect 5935 -515 6000 -500
rect 5950 -550 6000 -515
rect 6100 -535 6150 -450
rect 6400 -500 6650 -450
rect 6100 -550 6165 -535
rect 4900 -600 5150 -550
rect 5400 -600 5650 -550
rect 5750 -600 5900 -550
rect 5985 -565 6050 -550
rect 6000 -600 6050 -565
rect 6150 -600 6350 -550
rect 6400 -600 6450 -500
rect 6600 -600 6650 -500
rect 6750 -550 6800 -350
rect 6835 -365 6965 -350
rect 6850 -400 6950 -365
rect 6890 -410 6910 -400
rect 7000 -550 7050 -350
rect 7150 -315 7215 -300
rect 7385 -315 7450 -300
rect 7150 -385 7200 -315
rect 7400 -350 7450 -315
rect 7150 -400 7215 -385
rect 7200 -450 7400 -400
rect 7385 -465 7450 -450
rect 7150 -535 7200 -500
rect 7400 -535 7450 -465
rect 7150 -550 7215 -535
rect 7385 -550 7450 -535
rect 6700 -600 6850 -550
rect 6950 -600 7100 -550
rect 7200 -600 7400 -550
rect -1000 -800 -750 -750
rect -650 -800 -600 -750
rect -350 -800 -300 -750
rect -950 -900 -900 -800
rect -765 -815 -700 -800
rect -615 -815 -550 -800
rect -750 -885 -700 -815
rect -765 -900 -700 -885
rect -600 -900 -550 -815
rect -400 -815 -335 -800
rect -400 -900 -350 -815
rect -200 -900 -150 -850
rect -950 -950 -750 -900
rect -565 -915 -500 -900
rect -550 -950 -500 -915
rect -450 -915 -385 -900
rect -450 -950 -400 -915
rect -950 -1050 -900 -950
rect -765 -965 -700 -950
rect -515 -965 -435 -950
rect -750 -1035 -700 -965
rect -765 -1050 -700 -1035
rect -500 -1050 -450 -965
rect -200 -1000 -150 -950
rect -1000 -1100 -750 -1050
rect -550 -1100 -400 -1050
rect -950 -1300 -750 -1250
rect -1000 -1315 -935 -1300
rect -765 -1315 -700 -1300
rect -1000 -1385 -950 -1315
rect -750 -1350 -700 -1315
rect -1000 -1400 -935 -1385
rect -950 -1450 -750 -1400
rect -765 -1465 -700 -1450
rect -1000 -1535 -950 -1500
rect -750 -1535 -700 -1465
rect -1000 -1550 -935 -1535
rect -765 -1550 -700 -1535
rect -650 -1535 -600 -1250
rect -450 -1500 -400 -1250
rect -300 -1300 -100 -1250
rect 150 -1285 200 -1250
rect 149 -1300 201 -1285
rect 350 -1300 600 -1250
rect 750 -1300 950 -1250
rect 1050 -1300 1200 -1250
rect 1250 -1300 1400 -1250
rect 1550 -1285 1600 -1250
rect 1549 -1300 1601 -1285
rect 1750 -1300 1800 -1250
rect 2000 -1300 2100 -1250
rect 2250 -1285 2300 -1250
rect 2249 -1300 2301 -1285
rect 2600 -1300 2750 -1250
rect 2850 -1285 2950 -1250
rect 2835 -1300 2950 -1285
rect 3200 -1300 3400 -1250
rect -500 -1535 -400 -1500
rect -650 -1550 -585 -1535
rect -515 -1550 -400 -1535
rect -250 -1550 -200 -1300
rect -115 -1315 -50 -1300
rect -100 -1350 -50 -1315
rect 100 -1315 164 -1300
rect 186 -1315 250 -1300
rect 100 -1350 150 -1315
rect 200 -1350 250 -1315
rect -65 -1365 0 -1350
rect -50 -1535 0 -1365
rect -65 -1550 0 -1535
rect 50 -1365 115 -1350
rect 235 -1365 300 -1350
rect 50 -1450 100 -1365
rect 250 -1450 300 -1365
rect 50 -1500 300 -1450
rect -950 -1600 -750 -1550
rect -600 -1600 -500 -1550
rect -450 -1600 -350 -1550
rect -300 -1600 -50 -1550
rect 50 -1600 100 -1500
rect 250 -1600 300 -1500
rect 400 -1400 450 -1300
rect 585 -1315 650 -1300
rect 600 -1385 650 -1315
rect 585 -1400 650 -1385
rect 700 -1315 765 -1300
rect 935 -1315 1000 -1300
rect 700 -1385 750 -1315
rect 950 -1350 1000 -1315
rect 700 -1400 765 -1385
rect 1100 -1400 1150 -1300
rect 1300 -1400 1350 -1300
rect 1500 -1315 1564 -1300
rect 1586 -1315 1650 -1300
rect 1785 -1315 1850 -1300
rect 1500 -1350 1550 -1315
rect 1600 -1350 1650 -1315
rect 1800 -1350 1850 -1315
rect 400 -1450 600 -1400
rect 750 -1450 950 -1400
rect 1100 -1450 1350 -1400
rect 400 -1550 450 -1450
rect 500 -1500 550 -1450
rect 935 -1465 1000 -1450
rect 535 -1515 600 -1500
rect 550 -1550 600 -1515
rect 700 -1535 750 -1500
rect 950 -1535 1000 -1465
rect 700 -1550 765 -1535
rect 935 -1550 1000 -1535
rect 1100 -1550 1150 -1450
rect 1300 -1550 1350 -1450
rect 1450 -1365 1515 -1350
rect 1635 -1365 1700 -1350
rect 1450 -1450 1500 -1365
rect 1650 -1450 1700 -1365
rect 1450 -1500 1700 -1450
rect 350 -1600 500 -1550
rect 585 -1565 650 -1550
rect 600 -1600 650 -1565
rect 750 -1600 950 -1550
rect 1050 -1600 1200 -1550
rect 1250 -1600 1400 -1550
rect 1450 -1600 1500 -1500
rect 1650 -1600 1700 -1500
rect 1800 -1400 1900 -1350
rect 1800 -1550 1850 -1400
rect 1885 -1415 1950 -1400
rect 1900 -1450 1950 -1415
rect 2000 -1450 2050 -1300
rect 2200 -1315 2264 -1300
rect 2286 -1315 2350 -1300
rect 2200 -1350 2250 -1315
rect 2300 -1350 2350 -1315
rect 1935 -1465 2050 -1450
rect 1950 -1500 2050 -1465
rect 1750 -1600 1900 -1550
rect 2000 -1600 2050 -1500
rect 2150 -1365 2215 -1350
rect 2335 -1365 2400 -1350
rect 2150 -1450 2200 -1365
rect 2350 -1450 2400 -1365
rect 2150 -1500 2400 -1450
rect 2150 -1600 2200 -1500
rect 2350 -1600 2400 -1500
rect 2650 -1400 2700 -1300
rect 2800 -1385 2850 -1300
rect 2785 -1400 2850 -1385
rect 3150 -1315 3215 -1300
rect 3385 -1315 3450 -1300
rect 3150 -1385 3200 -1315
rect 3400 -1350 3450 -1315
rect 3150 -1400 3215 -1385
rect 2650 -1450 2800 -1400
rect 3200 -1450 3400 -1400
rect 2650 -1550 2700 -1450
rect 2785 -1465 2850 -1450
rect 3385 -1465 3450 -1450
rect 2800 -1550 2850 -1465
rect 3150 -1535 3200 -1500
rect 3400 -1535 3450 -1465
rect 3150 -1550 3215 -1535
rect 3385 -1550 3450 -1535
rect 2500 -1600 2550 -1550
rect 2600 -1600 2750 -1550
rect 2835 -1565 2950 -1550
rect 2850 -1600 2950 -1565
rect 3050 -1600 3100 -1550
rect 3200 -1600 3400 -1550
rect -1000 -1785 -950 -1750
rect -700 -1785 -650 -1750
rect -1000 -1800 -935 -1785
rect -715 -1800 -650 -1785
rect -600 -1800 -450 -1750
rect -400 -1800 -150 -1750
rect 50 -1785 100 -1750
rect 49 -1800 101 -1785
rect 350 -1800 550 -1750
rect 750 -1800 1000 -1750
rect 1100 -1800 1250 -1750
rect 1300 -1800 1450 -1750
rect 1600 -1785 1650 -1750
rect 1599 -1800 1651 -1785
rect 1850 -1800 2100 -1750
rect 2350 -1800 2600 -1750
rect -950 -1935 -900 -1800
rect -750 -1935 -700 -1800
rect -950 -1950 -885 -1935
rect -765 -1950 -700 -1935
rect -900 -2035 -850 -1950
rect -800 -2035 -750 -1950
rect -900 -2050 -836 -2035
rect -814 -2050 -750 -2035
rect -550 -2050 -500 -1800
rect -350 -1900 -300 -1800
rect -165 -1815 -100 -1800
rect -150 -1885 -100 -1815
rect 0 -1815 64 -1800
rect 86 -1815 150 -1800
rect 0 -1850 50 -1815
rect 100 -1850 150 -1815
rect -165 -1900 -100 -1885
rect -50 -1865 15 -1850
rect 135 -1865 200 -1850
rect -350 -1950 -150 -1900
rect -50 -1950 0 -1865
rect 150 -1950 200 -1865
rect -350 -2050 -300 -1950
rect -250 -2000 -200 -1950
rect -50 -2000 200 -1950
rect -215 -2015 -150 -2000
rect -200 -2050 -150 -2015
rect -851 -2065 -799 -2050
rect -850 -2100 -800 -2065
rect -600 -2100 -450 -2050
rect -400 -2100 -250 -2050
rect -165 -2065 -100 -2050
rect -150 -2100 -100 -2065
rect -50 -2100 0 -2000
rect 150 -2100 200 -2000
rect 250 -2035 300 -2000
rect 450 -2035 500 -1800
rect 250 -2050 315 -2035
rect 435 -2050 500 -2035
rect 800 -1900 850 -1800
rect 985 -1815 1050 -1800
rect 1000 -1885 1050 -1815
rect 985 -1900 1050 -1885
rect 1150 -1900 1200 -1800
rect 1350 -1900 1400 -1800
rect 1550 -1815 1614 -1800
rect 1636 -1815 1700 -1800
rect 1550 -1850 1600 -1815
rect 1650 -1850 1700 -1815
rect 1800 -1815 1865 -1800
rect 1800 -1850 1850 -1815
rect 800 -1950 1000 -1900
rect 1150 -1950 1400 -1900
rect 800 -2050 850 -1950
rect 985 -1965 1050 -1950
rect 1000 -2035 1050 -1965
rect 985 -2050 1050 -2035
rect 1150 -2050 1200 -1950
rect 1350 -2050 1400 -1950
rect 1500 -1865 1565 -1850
rect 1685 -1865 1750 -1850
rect 1500 -1950 1550 -1865
rect 1700 -1950 1750 -1865
rect 1500 -2000 1750 -1950
rect 300 -2100 450 -2050
rect 750 -2100 1000 -2050
rect 1100 -2100 1250 -2050
rect 1300 -2100 1450 -2050
rect 1500 -2100 1550 -2000
rect 1700 -2100 1750 -2000
rect 1950 -2050 2000 -1800
rect 2085 -1815 2150 -1800
rect 2100 -1850 2150 -1815
rect 2400 -1900 2450 -1800
rect 2585 -1815 2650 -1800
rect 2600 -1885 2650 -1815
rect 2585 -1900 2650 -1885
rect 2400 -1950 2600 -1900
rect 2400 -2050 2450 -1950
rect 2585 -1965 2650 -1950
rect 2600 -2035 2650 -1965
rect 2585 -2050 2650 -2035
rect 1900 -2100 2050 -2050
rect 2250 -2100 2300 -2050
rect 2350 -2100 2600 -2050
rect -950 -2300 -750 -2250
rect -650 -2300 -500 -2250
rect -450 -2300 -300 -2250
rect -250 -2300 0 -2250
rect 150 -2300 350 -2250
rect 400 -2300 450 -2250
rect 700 -2300 750 -2250
rect 900 -2285 950 -2250
rect 899 -2300 951 -2285
rect 1150 -2300 1350 -2250
rect 1650 -2300 1800 -2250
rect 1950 -2300 2100 -2250
rect 2200 -2300 2350 -2250
rect 2500 -2300 2650 -2250
rect 2700 -2300 2900 -2250
rect 3150 -2285 3200 -2250
rect 3149 -2300 3201 -2285
rect 3500 -2300 3750 -2250
rect 4000 -2300 4050 -2250
rect 4250 -2300 4350 -2250
rect -1000 -2315 -935 -2300
rect -765 -2315 -700 -2300
rect -1000 -2385 -950 -2315
rect -750 -2350 -700 -2315
rect -1000 -2400 -935 -2385
rect -600 -2400 -550 -2300
rect -400 -2400 -350 -2300
rect -950 -2450 -750 -2400
rect -600 -2450 -350 -2400
rect -765 -2465 -700 -2450
rect -1000 -2535 -950 -2500
rect -750 -2535 -700 -2465
rect -1000 -2550 -935 -2535
rect -765 -2550 -700 -2535
rect -600 -2550 -550 -2450
rect -400 -2550 -350 -2450
rect -200 -2400 -150 -2300
rect -15 -2315 50 -2300
rect 0 -2385 50 -2315
rect -15 -2400 50 -2385
rect 100 -2315 165 -2300
rect 435 -2315 500 -2300
rect 100 -2400 150 -2315
rect 450 -2400 500 -2315
rect 650 -2315 715 -2300
rect 850 -2315 914 -2300
rect 936 -2315 1000 -2300
rect 650 -2400 700 -2315
rect 850 -2350 900 -2315
rect 950 -2350 1000 -2315
rect 1100 -2315 1165 -2300
rect 1335 -2315 1400 -2300
rect 800 -2365 865 -2350
rect 985 -2365 1050 -2350
rect -200 -2450 0 -2400
rect 100 -2450 300 -2400
rect 485 -2415 550 -2400
rect 500 -2450 550 -2415
rect 600 -2415 665 -2400
rect 600 -2450 650 -2415
rect 800 -2450 850 -2365
rect 1000 -2450 1050 -2365
rect 1100 -2385 1150 -2315
rect 1350 -2350 1400 -2315
rect 1600 -2315 1665 -2300
rect 1785 -2315 1850 -2300
rect 1100 -2400 1165 -2385
rect 1150 -2450 1350 -2400
rect -200 -2550 -150 -2450
rect -100 -2500 -50 -2450
rect -65 -2515 0 -2500
rect -50 -2550 0 -2515
rect 100 -2535 150 -2450
rect 535 -2465 615 -2450
rect 100 -2550 165 -2535
rect 550 -2550 600 -2465
rect 800 -2500 1050 -2450
rect 1335 -2465 1400 -2450
rect -950 -2600 -750 -2550
rect -650 -2600 -500 -2550
rect -450 -2600 -300 -2550
rect -250 -2600 -100 -2550
rect -15 -2565 50 -2550
rect 0 -2600 50 -2565
rect 150 -2600 350 -2550
rect 500 -2600 650 -2550
rect 800 -2600 850 -2500
rect 1000 -2600 1050 -2500
rect 1100 -2535 1150 -2500
rect 1350 -2535 1400 -2465
rect 1100 -2550 1165 -2535
rect 1335 -2550 1400 -2535
rect 1600 -2535 1650 -2315
rect 1800 -2350 1850 -2315
rect 1900 -2315 1965 -2300
rect 2085 -2315 2150 -2300
rect 1750 -2500 1850 -2450
rect 1800 -2535 1850 -2500
rect 1600 -2550 1665 -2535
rect 1785 -2550 1850 -2535
rect 1900 -2535 1950 -2315
rect 2100 -2535 2150 -2315
rect 2250 -2485 2300 -2300
rect 2250 -2500 2315 -2485
rect 1900 -2550 1965 -2535
rect 2085 -2550 2150 -2535
rect 2300 -2535 2350 -2500
rect 2400 -2535 2450 -2450
rect 2550 -2485 2600 -2300
rect 2535 -2500 2600 -2485
rect 2500 -2535 2550 -2500
rect 2300 -2550 2364 -2535
rect 2386 -2550 2464 -2535
rect 2486 -2550 2550 -2535
rect 2750 -2550 2800 -2300
rect 2885 -2315 2950 -2300
rect 2900 -2350 2950 -2315
rect 3100 -2315 3164 -2300
rect 3186 -2315 3250 -2300
rect 3100 -2350 3150 -2315
rect 3200 -2350 3250 -2315
rect 2935 -2365 3000 -2350
rect 2950 -2535 3000 -2365
rect 2935 -2550 3000 -2535
rect 3050 -2365 3115 -2350
rect 3235 -2365 3300 -2350
rect 3050 -2450 3100 -2365
rect 3250 -2450 3300 -2365
rect 3050 -2500 3300 -2450
rect 1150 -2600 1350 -2550
rect 1650 -2600 1800 -2550
rect 1950 -2600 2100 -2550
rect 2349 -2565 2401 -2550
rect 2449 -2565 2501 -2550
rect 2350 -2600 2400 -2565
rect 2450 -2600 2500 -2565
rect 2700 -2600 2950 -2550
rect 3050 -2600 3100 -2500
rect 3250 -2600 3300 -2500
rect 3550 -2400 3600 -2300
rect 3735 -2315 3800 -2300
rect 4035 -2315 4100 -2300
rect 3750 -2385 3800 -2315
rect 3735 -2400 3800 -2385
rect 4050 -2350 4100 -2315
rect 4050 -2400 4150 -2350
rect 3550 -2450 3750 -2400
rect 3550 -2550 3600 -2450
rect 3735 -2465 3800 -2450
rect 3750 -2535 3800 -2465
rect 3735 -2550 3800 -2535
rect 4050 -2550 4100 -2400
rect 4135 -2415 4200 -2400
rect 4150 -2450 4200 -2415
rect 4250 -2450 4300 -2300
rect 4185 -2465 4300 -2450
rect 4200 -2500 4300 -2465
rect 3400 -2600 3450 -2550
rect 3500 -2600 3750 -2550
rect 3900 -2600 3950 -2550
rect 4000 -2600 4150 -2550
rect 4250 -2600 4300 -2500
rect -950 -2800 -750 -2750
rect -1000 -2815 -935 -2800
rect -765 -2815 -700 -2800
rect -1000 -2885 -950 -2815
rect -750 -2850 -700 -2815
rect -1000 -2900 -935 -2885
rect -950 -2950 -750 -2900
rect -765 -2965 -700 -2950
rect -1000 -3035 -950 -3000
rect -750 -3035 -700 -2965
rect -1000 -3050 -935 -3035
rect -765 -3050 -700 -3035
rect -650 -3035 -600 -2750
rect -450 -3000 -400 -2750
rect -300 -2800 -100 -2750
rect 50 -2800 200 -2750
rect 250 -2800 400 -2750
rect 550 -2785 600 -2750
rect 549 -2800 601 -2785
rect 750 -2800 1000 -2750
rect 1150 -2800 1350 -2750
rect 1550 -2785 1600 -2750
rect 1549 -2800 1601 -2785
rect 1750 -2800 1800 -2750
rect 2000 -2800 2100 -2750
rect 2350 -2800 2550 -2750
rect -500 -3035 -400 -3000
rect -650 -3050 -585 -3035
rect -515 -3050 -400 -3035
rect -250 -3050 -200 -2800
rect -115 -2815 -50 -2800
rect -100 -2850 -50 -2815
rect -65 -2865 0 -2850
rect -50 -3035 0 -2865
rect -65 -3050 0 -3035
rect 100 -2900 150 -2800
rect 300 -2900 350 -2800
rect 500 -2815 564 -2800
rect 586 -2815 650 -2800
rect 500 -2850 550 -2815
rect 600 -2850 650 -2815
rect 100 -2950 350 -2900
rect 100 -3050 150 -2950
rect 300 -3050 350 -2950
rect 450 -2865 515 -2850
rect 635 -2865 700 -2850
rect 450 -2950 500 -2865
rect 650 -2950 700 -2865
rect 450 -3000 700 -2950
rect -950 -3100 -750 -3050
rect -600 -3100 -500 -3050
rect -450 -3100 -350 -3050
rect -300 -3100 -50 -3050
rect 50 -3100 200 -3050
rect 250 -3100 400 -3050
rect 450 -3100 500 -3000
rect 650 -3100 700 -3000
rect 800 -2900 850 -2800
rect 985 -2815 1050 -2800
rect 1000 -2885 1050 -2815
rect 985 -2900 1050 -2885
rect 1100 -2815 1165 -2800
rect 1335 -2815 1400 -2800
rect 1100 -2885 1150 -2815
rect 1350 -2850 1400 -2815
rect 1500 -2815 1564 -2800
rect 1586 -2815 1650 -2800
rect 1785 -2815 1850 -2800
rect 1500 -2850 1550 -2815
rect 1600 -2850 1650 -2815
rect 1800 -2850 1850 -2815
rect 1450 -2865 1515 -2850
rect 1635 -2865 1700 -2850
rect 1100 -2900 1165 -2885
rect 800 -2950 1000 -2900
rect 1150 -2950 1350 -2900
rect 1450 -2950 1500 -2865
rect 1650 -2950 1700 -2865
rect 800 -3050 850 -2950
rect 900 -3000 950 -2950
rect 1335 -2965 1400 -2950
rect 935 -3015 1000 -3000
rect 950 -3050 1000 -3015
rect 1100 -3035 1150 -3000
rect 1350 -3035 1400 -2965
rect 1100 -3050 1165 -3035
rect 1335 -3050 1400 -3035
rect 1450 -3000 1700 -2950
rect 750 -3100 900 -3050
rect 985 -3065 1050 -3050
rect 1000 -3100 1050 -3065
rect 1150 -3100 1350 -3050
rect 1450 -3100 1500 -3000
rect 1650 -3100 1700 -3000
rect 1800 -2900 1900 -2850
rect 1800 -3050 1850 -2900
rect 1885 -2915 1950 -2900
rect 1900 -2950 1950 -2915
rect 2000 -2950 2050 -2800
rect 2300 -2815 2365 -2800
rect 2535 -2815 2600 -2800
rect 2300 -2885 2350 -2815
rect 2550 -2850 2600 -2815
rect 2300 -2900 2365 -2885
rect 2350 -2950 2550 -2900
rect 1935 -2965 2050 -2950
rect 2535 -2965 2600 -2950
rect 1950 -3000 2050 -2965
rect 1750 -3100 1900 -3050
rect 2000 -3100 2050 -3000
rect 2300 -3035 2350 -3000
rect 2550 -3035 2600 -2965
rect 2300 -3050 2365 -3035
rect 2535 -3050 2600 -3035
rect 2200 -3100 2250 -3050
rect 2350 -3100 2550 -3050
<< end >>
