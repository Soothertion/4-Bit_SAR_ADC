** sch_path: /home/ttuser/Desktop/NComp.sch
.subckt NComp VPWR Vref Vin Vcomp_n VGND
*.PININFO Vcomp_n:O Vin:I Vref:I VPWR:I VGND:I
XM29 VGND Vref net4 VGND sky130_fd_pr__nfet_01v8_lvt L=4 W=2 nf=1 m=1
XM30 VGND Vin net3 VGND sky130_fd_pr__nfet_01v8_lvt L=4 W=2 nf=1 m=1
XM31 VPWR net4 net4 VPWR sky130_fd_pr__pfet_01v8_lvt L=1 W=4 nf=1 m=1
XM32 VPWR net3 net3 VPWR sky130_fd_pr__pfet_01v8_lvt L=1 W=4 nf=1 m=1
XM33 VPWR net3 net1 VPWR sky130_fd_pr__pfet_01v8_lvt L=2 W=4 nf=1 m=1
XM34 VPWR net4 net2 VPWR sky130_fd_pr__pfet_01v8_lvt L=2 W=4 nf=1 m=1
XM35 VGND net2 net2 VGND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=2 m=1
XM36 VGND net2 net1 VGND sky130_fd_pr__nfet_01v8_lvt L=2 W=8 nf=2 m=1
XM37 Vcomp_n net1 VPWR VPWR sky130_fd_pr__pfet_01v8_lvt L=0.5 W=0.5 nf=1 m=1
XM38 Vcomp_n net1 VGND VGND sky130_fd_pr__nfet_01v8_lvt L=0.5 W=1.8 nf=1 m=1
.ends
.end
