** sch_path: /home/ttuser/Desktop/DAC.sch
.subckt DAC Vdac D0 D2 D3 D1 VGND
*.PININFO Vdac:O D0:I D1:I D2:I D3:I VGND:I
XR1 VGND net1 VGND sky130_fd_pr__res_high_po_0p35 L=12 mult=1 m=1
XR9 net1 net2 VGND sky130_fd_pr__res_high_po_0p35 L=4.8 mult=1 m=1
XR2 net2 net3 VGND sky130_fd_pr__res_high_po_0p35 L=4.8 mult=1 m=1
XR3 net3 Vdac VGND sky130_fd_pr__res_high_po_0p35 L=4.8 mult=1 m=1
XR4 D0 net1 VGND sky130_fd_pr__res_high_po_0p35 L=10.2 mult=1 m=1
XR5 D1 net2 VGND sky130_fd_pr__res_high_po_0p35 L=9.8 mult=1 m=1
XR6 D2 net3 VGND sky130_fd_pr__res_high_po_0p35 L=9.8 mult=1 m=1
XR7 D3 Vdac VGND sky130_fd_pr__res_high_po_0p35 L=10 mult=1 m=1
.ends
.end
