magic
tech sky130A
magscale 1 2
timestamp 1740303368
<< viali >>
rect 1409 7497 1443 7531
rect 1593 7361 1627 7395
rect 1869 7361 1903 7395
rect 2053 7361 2087 7395
rect 1685 7157 1719 7191
rect 2237 7157 2271 7191
rect 4905 6681 4939 6715
rect 6193 6613 6227 6647
rect 4353 6273 4387 6307
rect 2513 6205 2547 6239
rect 2881 6205 2915 6239
rect 4813 6069 4847 6103
rect 3801 5865 3835 5899
rect 4123 5865 4157 5899
rect 1869 5729 1903 5763
rect 3295 5729 3329 5763
rect 5549 5729 5583 5763
rect 5825 5729 5859 5763
rect 1593 5661 1627 5695
rect 3617 5593 3651 5627
rect 3157 5321 3191 5355
rect 1593 5185 1627 5219
rect 3617 5185 3651 5219
rect 5457 5185 5491 5219
rect 6653 5185 6687 5219
rect 5089 5117 5123 5151
rect 6469 5049 6503 5083
rect 1409 4981 1443 5015
rect 1869 4641 1903 4675
rect 5733 4641 5767 4675
rect 6101 4641 6135 4675
rect 1593 4573 1627 4607
rect 3295 4573 3329 4607
rect 4261 4573 4295 4607
rect 3617 4505 3651 4539
rect 3801 4437 3835 4471
rect 2329 4233 2363 4267
rect 2789 4097 2823 4131
rect 4261 4097 4295 4131
rect 4629 4097 4663 4131
rect 3893 3689 3927 3723
rect 3295 3621 3329 3655
rect 1869 3553 1903 3587
rect 5457 3553 5491 3587
rect 5825 3553 5859 3587
rect 1593 3485 1627 3519
rect 3617 3485 3651 3519
rect 4169 3349 4203 3383
rect 1593 3009 1627 3043
rect 1869 3009 1903 3043
rect 2605 3009 2639 3043
rect 4077 3009 4111 3043
rect 2145 2941 2179 2975
rect 4445 2941 4479 2975
rect 1409 2873 1443 2907
rect 1685 2805 1719 2839
rect 1685 2601 1719 2635
rect 3433 2601 3467 2635
rect 4261 2601 4295 2635
rect 3157 2397 3191 2431
rect 3617 2397 3651 2431
rect 5549 2397 5583 2431
<< metal1 >>
rect 1104 7642 6992 7664
rect 1104 7590 2658 7642
rect 2710 7590 2722 7642
rect 2774 7590 2786 7642
rect 2838 7590 2850 7642
rect 2902 7590 2914 7642
rect 2966 7590 2978 7642
rect 3030 7590 4158 7642
rect 4210 7590 4222 7642
rect 4274 7590 4286 7642
rect 4338 7590 4350 7642
rect 4402 7590 4414 7642
rect 4466 7590 4478 7642
rect 4530 7590 5658 7642
rect 5710 7590 5722 7642
rect 5774 7590 5786 7642
rect 5838 7590 5850 7642
rect 5902 7590 5914 7642
rect 5966 7590 5978 7642
rect 6030 7590 6992 7642
rect 1104 7568 6992 7590
rect 1394 7488 1400 7540
rect 1452 7488 1458 7540
rect 1581 7395 1639 7401
rect 1581 7361 1593 7395
rect 1627 7361 1639 7395
rect 1581 7355 1639 7361
rect 1857 7395 1915 7401
rect 1857 7361 1869 7395
rect 1903 7361 1915 7395
rect 1857 7355 1915 7361
rect 1596 7256 1624 7355
rect 1872 7324 1900 7355
rect 2038 7352 2044 7404
rect 2096 7352 2102 7404
rect 3142 7324 3148 7336
rect 1872 7296 3148 7324
rect 3142 7284 3148 7296
rect 3200 7284 3206 7336
rect 4062 7256 4068 7268
rect 1596 7228 4068 7256
rect 4062 7216 4068 7228
rect 4120 7216 4126 7268
rect 1670 7148 1676 7200
rect 1728 7148 1734 7200
rect 2225 7191 2283 7197
rect 2225 7157 2237 7191
rect 2271 7188 2283 7191
rect 3050 7188 3056 7200
rect 2271 7160 3056 7188
rect 2271 7157 2283 7160
rect 2225 7151 2283 7157
rect 3050 7148 3056 7160
rect 3108 7148 3114 7200
rect 1104 7098 6992 7120
rect 1104 7046 1918 7098
rect 1970 7046 1982 7098
rect 2034 7046 2046 7098
rect 2098 7046 2110 7098
rect 2162 7046 2174 7098
rect 2226 7046 2238 7098
rect 2290 7046 3418 7098
rect 3470 7046 3482 7098
rect 3534 7046 3546 7098
rect 3598 7046 3610 7098
rect 3662 7046 3674 7098
rect 3726 7046 3738 7098
rect 3790 7046 4918 7098
rect 4970 7046 4982 7098
rect 5034 7046 5046 7098
rect 5098 7046 5110 7098
rect 5162 7046 5174 7098
rect 5226 7046 5238 7098
rect 5290 7046 6418 7098
rect 6470 7046 6482 7098
rect 6534 7046 6546 7098
rect 6598 7046 6610 7098
rect 6662 7046 6674 7098
rect 6726 7046 6738 7098
rect 6790 7046 6992 7098
rect 1104 7024 6992 7046
rect 4706 6672 4712 6724
rect 4764 6712 4770 6724
rect 4893 6715 4951 6721
rect 4893 6712 4905 6715
rect 4764 6684 4905 6712
rect 4764 6672 4770 6684
rect 4893 6681 4905 6684
rect 4939 6681 4951 6715
rect 4893 6675 4951 6681
rect 6178 6604 6184 6656
rect 6236 6604 6242 6656
rect 1104 6554 6992 6576
rect 1104 6502 2658 6554
rect 2710 6502 2722 6554
rect 2774 6502 2786 6554
rect 2838 6502 2850 6554
rect 2902 6502 2914 6554
rect 2966 6502 2978 6554
rect 3030 6502 4158 6554
rect 4210 6502 4222 6554
rect 4274 6502 4286 6554
rect 4338 6502 4350 6554
rect 4402 6502 4414 6554
rect 4466 6502 4478 6554
rect 4530 6502 5658 6554
rect 5710 6502 5722 6554
rect 5774 6502 5786 6554
rect 5838 6502 5850 6554
rect 5902 6502 5914 6554
rect 5966 6502 5978 6554
rect 6030 6502 6992 6554
rect 1104 6480 6992 6502
rect 3878 6332 3884 6384
rect 3936 6332 3942 6384
rect 4341 6307 4399 6313
rect 4341 6273 4353 6307
rect 4387 6273 4399 6307
rect 4341 6267 4399 6273
rect 2501 6239 2559 6245
rect 2501 6205 2513 6239
rect 2547 6236 2559 6239
rect 2866 6236 2872 6248
rect 2547 6208 2872 6236
rect 2547 6205 2559 6208
rect 2501 6199 2559 6205
rect 2866 6196 2872 6208
rect 2924 6196 2930 6248
rect 3970 6128 3976 6180
rect 4028 6168 4034 6180
rect 4356 6168 4384 6267
rect 4028 6140 4384 6168
rect 4028 6128 4034 6140
rect 4801 6103 4859 6109
rect 4801 6069 4813 6103
rect 4847 6100 4859 6103
rect 5442 6100 5448 6112
rect 4847 6072 5448 6100
rect 4847 6069 4859 6072
rect 4801 6063 4859 6069
rect 5442 6060 5448 6072
rect 5500 6060 5506 6112
rect 1104 6010 6992 6032
rect 1104 5958 1918 6010
rect 1970 5958 1982 6010
rect 2034 5958 2046 6010
rect 2098 5958 2110 6010
rect 2162 5958 2174 6010
rect 2226 5958 2238 6010
rect 2290 5958 3418 6010
rect 3470 5958 3482 6010
rect 3534 5958 3546 6010
rect 3598 5958 3610 6010
rect 3662 5958 3674 6010
rect 3726 5958 3738 6010
rect 3790 5958 4918 6010
rect 4970 5958 4982 6010
rect 5034 5958 5046 6010
rect 5098 5958 5110 6010
rect 5162 5958 5174 6010
rect 5226 5958 5238 6010
rect 5290 5958 6418 6010
rect 6470 5958 6482 6010
rect 6534 5958 6546 6010
rect 6598 5958 6610 6010
rect 6662 5958 6674 6010
rect 6726 5958 6738 6010
rect 6790 5958 6992 6010
rect 1104 5936 6992 5958
rect 3050 5856 3056 5908
rect 3108 5896 3114 5908
rect 3789 5899 3847 5905
rect 3108 5868 3188 5896
rect 3108 5856 3114 5868
rect 1857 5763 1915 5769
rect 1857 5729 1869 5763
rect 1903 5760 1915 5763
rect 3050 5760 3056 5772
rect 1903 5732 3056 5760
rect 1903 5729 1915 5732
rect 1857 5723 1915 5729
rect 3050 5720 3056 5732
rect 3108 5720 3114 5772
rect 1578 5652 1584 5704
rect 1636 5652 1642 5704
rect 3160 5624 3188 5868
rect 3789 5865 3801 5899
rect 3835 5896 3847 5899
rect 3878 5896 3884 5908
rect 3835 5868 3884 5896
rect 3835 5865 3847 5868
rect 3789 5859 3847 5865
rect 3878 5856 3884 5868
rect 3936 5856 3942 5908
rect 4062 5856 4068 5908
rect 4120 5905 4126 5908
rect 4120 5899 4169 5905
rect 4120 5865 4123 5899
rect 4157 5865 4169 5899
rect 4120 5859 4169 5865
rect 4120 5856 4126 5859
rect 3283 5763 3341 5769
rect 3283 5729 3295 5763
rect 3329 5760 3341 5763
rect 5537 5763 5595 5769
rect 5537 5760 5549 5763
rect 3329 5732 5549 5760
rect 3329 5729 3341 5732
rect 3283 5723 3341 5729
rect 5537 5729 5549 5732
rect 5583 5729 5595 5763
rect 5537 5723 5595 5729
rect 5813 5763 5871 5769
rect 5813 5729 5825 5763
rect 5859 5760 5871 5763
rect 6178 5760 6184 5772
rect 5859 5732 6184 5760
rect 5859 5729 5871 5732
rect 5813 5723 5871 5729
rect 6178 5720 6184 5732
rect 6236 5720 6242 5772
rect 3326 5624 3332 5636
rect 3082 5596 3332 5624
rect 3326 5584 3332 5596
rect 3384 5584 3390 5636
rect 3605 5627 3663 5633
rect 3605 5593 3617 5627
rect 3651 5624 3663 5627
rect 3970 5624 3976 5636
rect 3651 5596 3976 5624
rect 3651 5593 3663 5596
rect 3605 5587 3663 5593
rect 3970 5584 3976 5596
rect 4028 5584 4034 5636
rect 4062 5584 4068 5636
rect 4120 5624 4126 5636
rect 4120 5596 4370 5624
rect 4120 5584 4126 5596
rect 2866 5516 2872 5568
rect 2924 5556 2930 5568
rect 3878 5556 3884 5568
rect 2924 5528 3884 5556
rect 2924 5516 2930 5528
rect 3878 5516 3884 5528
rect 3936 5516 3942 5568
rect 1104 5466 6992 5488
rect 1104 5414 2658 5466
rect 2710 5414 2722 5466
rect 2774 5414 2786 5466
rect 2838 5414 2850 5466
rect 2902 5414 2914 5466
rect 2966 5414 2978 5466
rect 3030 5414 4158 5466
rect 4210 5414 4222 5466
rect 4274 5414 4286 5466
rect 4338 5414 4350 5466
rect 4402 5414 4414 5466
rect 4466 5414 4478 5466
rect 4530 5414 5658 5466
rect 5710 5414 5722 5466
rect 5774 5414 5786 5466
rect 5838 5414 5850 5466
rect 5902 5414 5914 5466
rect 5966 5414 5978 5466
rect 6030 5414 6992 5466
rect 1104 5392 6992 5414
rect 3142 5312 3148 5364
rect 3200 5312 3206 5364
rect 3976 5296 4028 5302
rect 3976 5238 4028 5244
rect 1581 5219 1639 5225
rect 1581 5185 1593 5219
rect 1627 5216 1639 5219
rect 2406 5216 2412 5228
rect 1627 5188 2412 5216
rect 1627 5185 1639 5188
rect 1581 5179 1639 5185
rect 2406 5176 2412 5188
rect 2464 5176 2470 5228
rect 3326 5176 3332 5228
rect 3384 5216 3390 5228
rect 3605 5219 3663 5225
rect 3605 5216 3617 5219
rect 3384 5188 3617 5216
rect 3384 5176 3390 5188
rect 3605 5185 3617 5188
rect 3651 5185 3663 5219
rect 3605 5179 3663 5185
rect 3620 5080 3648 5179
rect 5442 5176 5448 5228
rect 5500 5176 5506 5228
rect 6641 5219 6699 5225
rect 6641 5185 6653 5219
rect 6687 5216 6699 5219
rect 6914 5216 6920 5228
rect 6687 5188 6920 5216
rect 6687 5185 6699 5188
rect 6641 5179 6699 5185
rect 6914 5176 6920 5188
rect 6972 5176 6978 5228
rect 4614 5108 4620 5160
rect 4672 5148 4678 5160
rect 5077 5151 5135 5157
rect 5077 5148 5089 5151
rect 4672 5120 5089 5148
rect 4672 5108 4678 5120
rect 5077 5117 5089 5120
rect 5123 5148 5135 5151
rect 5123 5120 5488 5148
rect 5123 5117 5135 5120
rect 5077 5111 5135 5117
rect 5460 5092 5488 5120
rect 4062 5080 4068 5092
rect 3620 5052 4068 5080
rect 4062 5040 4068 5052
rect 4120 5040 4126 5092
rect 5442 5040 5448 5092
rect 5500 5080 5506 5092
rect 6457 5083 6515 5089
rect 6457 5080 6469 5083
rect 5500 5052 6469 5080
rect 5500 5040 5506 5052
rect 6457 5049 6469 5052
rect 6503 5049 6515 5083
rect 6457 5043 6515 5049
rect 842 4972 848 5024
rect 900 5012 906 5024
rect 1397 5015 1455 5021
rect 1397 5012 1409 5015
rect 900 4984 1409 5012
rect 900 4972 906 4984
rect 1397 4981 1409 4984
rect 1443 4981 1455 5015
rect 1397 4975 1455 4981
rect 1104 4922 6992 4944
rect 1104 4870 1918 4922
rect 1970 4870 1982 4922
rect 2034 4870 2046 4922
rect 2098 4870 2110 4922
rect 2162 4870 2174 4922
rect 2226 4870 2238 4922
rect 2290 4870 3418 4922
rect 3470 4870 3482 4922
rect 3534 4870 3546 4922
rect 3598 4870 3610 4922
rect 3662 4870 3674 4922
rect 3726 4870 3738 4922
rect 3790 4870 4918 4922
rect 4970 4870 4982 4922
rect 5034 4870 5046 4922
rect 5098 4870 5110 4922
rect 5162 4870 5174 4922
rect 5226 4870 5238 4922
rect 5290 4870 6418 4922
rect 6470 4870 6482 4922
rect 6534 4870 6546 4922
rect 6598 4870 6610 4922
rect 6662 4870 6674 4922
rect 6726 4870 6738 4922
rect 6790 4870 6992 4922
rect 1104 4848 6992 4870
rect 2406 4768 2412 4820
rect 2464 4808 2470 4820
rect 2464 4780 6132 4808
rect 2464 4768 2470 4780
rect 1857 4675 1915 4681
rect 1857 4641 1869 4675
rect 1903 4672 1915 4675
rect 3878 4672 3884 4684
rect 1903 4644 3884 4672
rect 1903 4641 1915 4644
rect 1857 4635 1915 4641
rect 3878 4632 3884 4644
rect 3936 4632 3942 4684
rect 5442 4632 5448 4684
rect 5500 4672 5506 4684
rect 6104 4681 6132 4780
rect 5721 4675 5779 4681
rect 5721 4672 5733 4675
rect 5500 4644 5733 4672
rect 5500 4632 5506 4644
rect 5721 4641 5733 4644
rect 5767 4641 5779 4675
rect 5721 4635 5779 4641
rect 6089 4675 6147 4681
rect 6089 4641 6101 4675
rect 6135 4641 6147 4675
rect 6089 4635 6147 4641
rect 1578 4564 1584 4616
rect 1636 4564 1642 4616
rect 3142 4564 3148 4616
rect 3200 4604 3206 4616
rect 3283 4607 3341 4613
rect 3283 4604 3295 4607
rect 3200 4576 3295 4604
rect 3200 4564 3206 4576
rect 3283 4573 3295 4576
rect 3329 4573 3341 4607
rect 3283 4567 3341 4573
rect 3786 4564 3792 4616
rect 3844 4604 3850 4616
rect 4062 4604 4068 4616
rect 3844 4576 4068 4604
rect 3844 4564 3850 4576
rect 4062 4564 4068 4576
rect 4120 4604 4126 4616
rect 4249 4607 4307 4613
rect 4249 4604 4261 4607
rect 4120 4576 4261 4604
rect 4120 4564 4126 4576
rect 4249 4573 4261 4576
rect 4295 4573 4307 4607
rect 4249 4567 4307 4573
rect 2498 4496 2504 4548
rect 2556 4496 2562 4548
rect 3605 4539 3663 4545
rect 3605 4505 3617 4539
rect 3651 4536 3663 4539
rect 3651 4508 4646 4536
rect 3651 4505 3663 4508
rect 3605 4499 3663 4505
rect 3789 4471 3847 4477
rect 3789 4437 3801 4471
rect 3835 4468 3847 4471
rect 4062 4468 4068 4480
rect 3835 4440 4068 4468
rect 3835 4437 3847 4440
rect 3789 4431 3847 4437
rect 4062 4428 4068 4440
rect 4120 4428 4126 4480
rect 1104 4378 6992 4400
rect 1104 4326 2658 4378
rect 2710 4326 2722 4378
rect 2774 4326 2786 4378
rect 2838 4326 2850 4378
rect 2902 4326 2914 4378
rect 2966 4326 2978 4378
rect 3030 4326 4158 4378
rect 4210 4326 4222 4378
rect 4274 4326 4286 4378
rect 4338 4326 4350 4378
rect 4402 4326 4414 4378
rect 4466 4326 4478 4378
rect 4530 4326 5658 4378
rect 5710 4326 5722 4378
rect 5774 4326 5786 4378
rect 5838 4326 5850 4378
rect 5902 4326 5914 4378
rect 5966 4326 5978 4378
rect 6030 4326 6992 4378
rect 1104 4304 6992 4326
rect 2317 4267 2375 4273
rect 2317 4233 2329 4267
rect 2363 4264 2375 4267
rect 2406 4264 2412 4276
rect 2363 4236 2412 4264
rect 2363 4233 2375 4236
rect 2317 4227 2375 4233
rect 2406 4224 2412 4236
rect 2464 4224 2470 4276
rect 3234 4224 3240 4276
rect 3292 4264 3298 4276
rect 3292 4236 4660 4264
rect 3292 4224 3298 4236
rect 3326 4156 3332 4208
rect 3384 4156 3390 4208
rect 2498 4088 2504 4140
rect 2556 4128 2562 4140
rect 2777 4131 2835 4137
rect 2777 4128 2789 4131
rect 2556 4100 2789 4128
rect 2556 4088 2562 4100
rect 2777 4097 2789 4100
rect 2823 4128 2835 4131
rect 3234 4128 3240 4140
rect 2823 4100 3240 4128
rect 2823 4097 2835 4100
rect 2777 4091 2835 4097
rect 3234 4088 3240 4100
rect 3292 4088 3298 4140
rect 4249 4131 4307 4137
rect 4249 4097 4261 4131
rect 4295 4128 4307 4131
rect 4522 4128 4528 4140
rect 4295 4100 4528 4128
rect 4295 4097 4307 4100
rect 4249 4091 4307 4097
rect 4522 4088 4528 4100
rect 4580 4088 4586 4140
rect 4632 4137 4660 4236
rect 4617 4131 4675 4137
rect 4617 4097 4629 4131
rect 4663 4097 4675 4131
rect 4617 4091 4675 4097
rect 3234 3884 3240 3936
rect 3292 3924 3298 3936
rect 3786 3924 3792 3936
rect 3292 3896 3792 3924
rect 3292 3884 3298 3896
rect 3786 3884 3792 3896
rect 3844 3884 3850 3936
rect 1104 3834 6992 3856
rect 1104 3782 1918 3834
rect 1970 3782 1982 3834
rect 2034 3782 2046 3834
rect 2098 3782 2110 3834
rect 2162 3782 2174 3834
rect 2226 3782 2238 3834
rect 2290 3782 3418 3834
rect 3470 3782 3482 3834
rect 3534 3782 3546 3834
rect 3598 3782 3610 3834
rect 3662 3782 3674 3834
rect 3726 3782 3738 3834
rect 3790 3782 4918 3834
rect 4970 3782 4982 3834
rect 5034 3782 5046 3834
rect 5098 3782 5110 3834
rect 5162 3782 5174 3834
rect 5226 3782 5238 3834
rect 5290 3782 6418 3834
rect 6470 3782 6482 3834
rect 6534 3782 6546 3834
rect 6598 3782 6610 3834
rect 6662 3782 6674 3834
rect 6726 3782 6738 3834
rect 6790 3782 6992 3834
rect 1104 3760 6992 3782
rect 3878 3680 3884 3732
rect 3936 3680 3942 3732
rect 3050 3612 3056 3664
rect 3108 3652 3114 3664
rect 3283 3655 3341 3661
rect 3283 3652 3295 3655
rect 3108 3624 3295 3652
rect 3108 3612 3114 3624
rect 3283 3621 3295 3624
rect 3329 3621 3341 3655
rect 3283 3615 3341 3621
rect 1857 3587 1915 3593
rect 1857 3553 1869 3587
rect 1903 3584 1915 3587
rect 3142 3584 3148 3596
rect 1903 3556 3148 3584
rect 1903 3553 1915 3556
rect 1857 3547 1915 3553
rect 3142 3544 3148 3556
rect 3200 3544 3206 3596
rect 3878 3544 3884 3596
rect 3936 3584 3942 3596
rect 5445 3587 5503 3593
rect 5445 3584 5457 3587
rect 3936 3556 5457 3584
rect 3936 3544 3942 3556
rect 5445 3553 5457 3556
rect 5491 3553 5503 3587
rect 5445 3547 5503 3553
rect 5813 3587 5871 3593
rect 5813 3553 5825 3587
rect 5859 3584 5871 3587
rect 6178 3584 6184 3596
rect 5859 3556 6184 3584
rect 5859 3553 5871 3556
rect 5813 3547 5871 3553
rect 6178 3544 6184 3556
rect 6236 3544 6242 3596
rect 1578 3476 1584 3528
rect 1636 3476 1642 3528
rect 3326 3476 3332 3528
rect 3384 3516 3390 3528
rect 3605 3519 3663 3525
rect 3605 3516 3617 3519
rect 3384 3488 3617 3516
rect 3384 3476 3390 3488
rect 3605 3485 3617 3488
rect 3651 3485 3663 3519
rect 3605 3479 3663 3485
rect 3234 3448 3240 3460
rect 3082 3420 3240 3448
rect 3234 3408 3240 3420
rect 3292 3448 3298 3460
rect 3292 3420 4462 3448
rect 3292 3408 3298 3420
rect 3970 3340 3976 3392
rect 4028 3380 4034 3392
rect 4157 3383 4215 3389
rect 4157 3380 4169 3383
rect 4028 3352 4169 3380
rect 4028 3340 4034 3352
rect 4157 3349 4169 3352
rect 4203 3349 4215 3383
rect 4157 3343 4215 3349
rect 1104 3290 6992 3312
rect 1104 3238 2658 3290
rect 2710 3238 2722 3290
rect 2774 3238 2786 3290
rect 2838 3238 2850 3290
rect 2902 3238 2914 3290
rect 2966 3238 2978 3290
rect 3030 3238 4158 3290
rect 4210 3238 4222 3290
rect 4274 3238 4286 3290
rect 4338 3238 4350 3290
rect 4402 3238 4414 3290
rect 4466 3238 4478 3290
rect 4530 3238 5658 3290
rect 5710 3238 5722 3290
rect 5774 3238 5786 3290
rect 5838 3238 5850 3290
rect 5902 3238 5914 3290
rect 5966 3238 5978 3290
rect 6030 3238 6992 3290
rect 1104 3216 6992 3238
rect 3970 3176 3976 3188
rect 3804 3148 3976 3176
rect 3804 3108 3832 3148
rect 3970 3136 3976 3148
rect 4028 3136 4034 3188
rect 3726 3080 3832 3108
rect 1581 3043 1639 3049
rect 1581 3009 1593 3043
rect 1627 3009 1639 3043
rect 1581 3003 1639 3009
rect 1857 3043 1915 3049
rect 1857 3009 1869 3043
rect 1903 3009 1915 3043
rect 1857 3003 1915 3009
rect 2593 3043 2651 3049
rect 2593 3009 2605 3043
rect 2639 3040 2651 3043
rect 3142 3040 3148 3052
rect 2639 3012 3148 3040
rect 2639 3009 2651 3012
rect 2593 3003 2651 3009
rect 842 2864 848 2916
rect 900 2904 906 2916
rect 1397 2907 1455 2913
rect 1397 2904 1409 2907
rect 900 2876 1409 2904
rect 900 2864 906 2876
rect 1397 2873 1409 2876
rect 1443 2873 1455 2907
rect 1596 2904 1624 3003
rect 1872 2972 1900 3003
rect 3142 3000 3148 3012
rect 3200 3000 3206 3052
rect 4065 3043 4123 3049
rect 4065 3009 4077 3043
rect 4111 3040 4123 3043
rect 4614 3040 4620 3052
rect 4111 3012 4620 3040
rect 4111 3009 4123 3012
rect 4065 3003 4123 3009
rect 4614 3000 4620 3012
rect 4672 3000 4678 3052
rect 2133 2975 2191 2981
rect 2133 2972 2145 2975
rect 1872 2944 2145 2972
rect 2133 2941 2145 2944
rect 2179 2941 2191 2975
rect 2133 2935 2191 2941
rect 4433 2975 4491 2981
rect 4433 2941 4445 2975
rect 4479 2941 4491 2975
rect 4433 2935 4491 2941
rect 1596 2876 3188 2904
rect 1397 2867 1455 2873
rect 1670 2796 1676 2848
rect 1728 2796 1734 2848
rect 3160 2836 3188 2876
rect 4062 2836 4068 2848
rect 3160 2808 4068 2836
rect 4062 2796 4068 2808
rect 4120 2836 4126 2848
rect 4448 2836 4476 2935
rect 4120 2808 4476 2836
rect 4120 2796 4126 2808
rect 1104 2746 6992 2768
rect 1104 2694 1918 2746
rect 1970 2694 1982 2746
rect 2034 2694 2046 2746
rect 2098 2694 2110 2746
rect 2162 2694 2174 2746
rect 2226 2694 2238 2746
rect 2290 2694 3418 2746
rect 3470 2694 3482 2746
rect 3534 2694 3546 2746
rect 3598 2694 3610 2746
rect 3662 2694 3674 2746
rect 3726 2694 3738 2746
rect 3790 2694 4918 2746
rect 4970 2694 4982 2746
rect 5034 2694 5046 2746
rect 5098 2694 5110 2746
rect 5162 2694 5174 2746
rect 5226 2694 5238 2746
rect 5290 2694 6418 2746
rect 6470 2694 6482 2746
rect 6534 2694 6546 2746
rect 6598 2694 6610 2746
rect 6662 2694 6674 2746
rect 6726 2694 6738 2746
rect 6790 2694 6992 2746
rect 1104 2672 6992 2694
rect 1578 2592 1584 2644
rect 1636 2632 1642 2644
rect 1673 2635 1731 2641
rect 1673 2632 1685 2635
rect 1636 2604 1685 2632
rect 1636 2592 1642 2604
rect 1673 2601 1685 2604
rect 1719 2601 1731 2635
rect 1673 2595 1731 2601
rect 3421 2635 3479 2641
rect 3421 2601 3433 2635
rect 3467 2632 3479 2635
rect 3878 2632 3884 2644
rect 3467 2604 3884 2632
rect 3467 2601 3479 2604
rect 3421 2595 3479 2601
rect 3878 2592 3884 2604
rect 3936 2592 3942 2644
rect 4249 2635 4307 2641
rect 4249 2601 4261 2635
rect 4295 2632 4307 2635
rect 4706 2632 4712 2644
rect 4295 2604 4712 2632
rect 4295 2601 4307 2604
rect 4249 2595 4307 2601
rect 4264 2496 4292 2595
rect 4706 2592 4712 2604
rect 4764 2592 4770 2644
rect 3160 2468 4292 2496
rect 3160 2437 3188 2468
rect 3145 2431 3203 2437
rect 3145 2397 3157 2431
rect 3191 2397 3203 2431
rect 3145 2391 3203 2397
rect 3605 2431 3663 2437
rect 3605 2397 3617 2431
rect 3651 2428 3663 2431
rect 3970 2428 3976 2440
rect 3651 2400 3976 2428
rect 3651 2397 3663 2400
rect 3605 2391 3663 2397
rect 3970 2388 3976 2400
rect 4028 2388 4034 2440
rect 5534 2388 5540 2440
rect 5592 2388 5598 2440
rect 1104 2202 6992 2224
rect 1104 2150 2658 2202
rect 2710 2150 2722 2202
rect 2774 2150 2786 2202
rect 2838 2150 2850 2202
rect 2902 2150 2914 2202
rect 2966 2150 2978 2202
rect 3030 2150 4158 2202
rect 4210 2150 4222 2202
rect 4274 2150 4286 2202
rect 4338 2150 4350 2202
rect 4402 2150 4414 2202
rect 4466 2150 4478 2202
rect 4530 2150 5658 2202
rect 5710 2150 5722 2202
rect 5774 2150 5786 2202
rect 5838 2150 5850 2202
rect 5902 2150 5914 2202
rect 5966 2150 5978 2202
rect 6030 2150 6992 2202
rect 1104 2128 6992 2150
<< via1 >>
rect 2658 7590 2710 7642
rect 2722 7590 2774 7642
rect 2786 7590 2838 7642
rect 2850 7590 2902 7642
rect 2914 7590 2966 7642
rect 2978 7590 3030 7642
rect 4158 7590 4210 7642
rect 4222 7590 4274 7642
rect 4286 7590 4338 7642
rect 4350 7590 4402 7642
rect 4414 7590 4466 7642
rect 4478 7590 4530 7642
rect 5658 7590 5710 7642
rect 5722 7590 5774 7642
rect 5786 7590 5838 7642
rect 5850 7590 5902 7642
rect 5914 7590 5966 7642
rect 5978 7590 6030 7642
rect 1400 7531 1452 7540
rect 1400 7497 1409 7531
rect 1409 7497 1443 7531
rect 1443 7497 1452 7531
rect 1400 7488 1452 7497
rect 2044 7395 2096 7404
rect 2044 7361 2053 7395
rect 2053 7361 2087 7395
rect 2087 7361 2096 7395
rect 2044 7352 2096 7361
rect 3148 7284 3200 7336
rect 4068 7216 4120 7268
rect 1676 7191 1728 7200
rect 1676 7157 1685 7191
rect 1685 7157 1719 7191
rect 1719 7157 1728 7191
rect 1676 7148 1728 7157
rect 3056 7148 3108 7200
rect 1918 7046 1970 7098
rect 1982 7046 2034 7098
rect 2046 7046 2098 7098
rect 2110 7046 2162 7098
rect 2174 7046 2226 7098
rect 2238 7046 2290 7098
rect 3418 7046 3470 7098
rect 3482 7046 3534 7098
rect 3546 7046 3598 7098
rect 3610 7046 3662 7098
rect 3674 7046 3726 7098
rect 3738 7046 3790 7098
rect 4918 7046 4970 7098
rect 4982 7046 5034 7098
rect 5046 7046 5098 7098
rect 5110 7046 5162 7098
rect 5174 7046 5226 7098
rect 5238 7046 5290 7098
rect 6418 7046 6470 7098
rect 6482 7046 6534 7098
rect 6546 7046 6598 7098
rect 6610 7046 6662 7098
rect 6674 7046 6726 7098
rect 6738 7046 6790 7098
rect 4712 6672 4764 6724
rect 6184 6647 6236 6656
rect 6184 6613 6193 6647
rect 6193 6613 6227 6647
rect 6227 6613 6236 6647
rect 6184 6604 6236 6613
rect 2658 6502 2710 6554
rect 2722 6502 2774 6554
rect 2786 6502 2838 6554
rect 2850 6502 2902 6554
rect 2914 6502 2966 6554
rect 2978 6502 3030 6554
rect 4158 6502 4210 6554
rect 4222 6502 4274 6554
rect 4286 6502 4338 6554
rect 4350 6502 4402 6554
rect 4414 6502 4466 6554
rect 4478 6502 4530 6554
rect 5658 6502 5710 6554
rect 5722 6502 5774 6554
rect 5786 6502 5838 6554
rect 5850 6502 5902 6554
rect 5914 6502 5966 6554
rect 5978 6502 6030 6554
rect 3884 6332 3936 6384
rect 2872 6239 2924 6248
rect 2872 6205 2881 6239
rect 2881 6205 2915 6239
rect 2915 6205 2924 6239
rect 2872 6196 2924 6205
rect 3976 6128 4028 6180
rect 5448 6060 5500 6112
rect 1918 5958 1970 6010
rect 1982 5958 2034 6010
rect 2046 5958 2098 6010
rect 2110 5958 2162 6010
rect 2174 5958 2226 6010
rect 2238 5958 2290 6010
rect 3418 5958 3470 6010
rect 3482 5958 3534 6010
rect 3546 5958 3598 6010
rect 3610 5958 3662 6010
rect 3674 5958 3726 6010
rect 3738 5958 3790 6010
rect 4918 5958 4970 6010
rect 4982 5958 5034 6010
rect 5046 5958 5098 6010
rect 5110 5958 5162 6010
rect 5174 5958 5226 6010
rect 5238 5958 5290 6010
rect 6418 5958 6470 6010
rect 6482 5958 6534 6010
rect 6546 5958 6598 6010
rect 6610 5958 6662 6010
rect 6674 5958 6726 6010
rect 6738 5958 6790 6010
rect 3056 5856 3108 5908
rect 3056 5720 3108 5772
rect 1584 5695 1636 5704
rect 1584 5661 1593 5695
rect 1593 5661 1627 5695
rect 1627 5661 1636 5695
rect 1584 5652 1636 5661
rect 3884 5856 3936 5908
rect 4068 5856 4120 5908
rect 6184 5720 6236 5772
rect 3332 5584 3384 5636
rect 3976 5584 4028 5636
rect 4068 5584 4120 5636
rect 2872 5516 2924 5568
rect 3884 5516 3936 5568
rect 2658 5414 2710 5466
rect 2722 5414 2774 5466
rect 2786 5414 2838 5466
rect 2850 5414 2902 5466
rect 2914 5414 2966 5466
rect 2978 5414 3030 5466
rect 4158 5414 4210 5466
rect 4222 5414 4274 5466
rect 4286 5414 4338 5466
rect 4350 5414 4402 5466
rect 4414 5414 4466 5466
rect 4478 5414 4530 5466
rect 5658 5414 5710 5466
rect 5722 5414 5774 5466
rect 5786 5414 5838 5466
rect 5850 5414 5902 5466
rect 5914 5414 5966 5466
rect 5978 5414 6030 5466
rect 3148 5355 3200 5364
rect 3148 5321 3157 5355
rect 3157 5321 3191 5355
rect 3191 5321 3200 5355
rect 3148 5312 3200 5321
rect 3976 5244 4028 5296
rect 2412 5176 2464 5228
rect 3332 5176 3384 5228
rect 5448 5219 5500 5228
rect 5448 5185 5457 5219
rect 5457 5185 5491 5219
rect 5491 5185 5500 5219
rect 5448 5176 5500 5185
rect 6920 5176 6972 5228
rect 4620 5108 4672 5160
rect 4068 5040 4120 5092
rect 5448 5040 5500 5092
rect 848 4972 900 5024
rect 1918 4870 1970 4922
rect 1982 4870 2034 4922
rect 2046 4870 2098 4922
rect 2110 4870 2162 4922
rect 2174 4870 2226 4922
rect 2238 4870 2290 4922
rect 3418 4870 3470 4922
rect 3482 4870 3534 4922
rect 3546 4870 3598 4922
rect 3610 4870 3662 4922
rect 3674 4870 3726 4922
rect 3738 4870 3790 4922
rect 4918 4870 4970 4922
rect 4982 4870 5034 4922
rect 5046 4870 5098 4922
rect 5110 4870 5162 4922
rect 5174 4870 5226 4922
rect 5238 4870 5290 4922
rect 6418 4870 6470 4922
rect 6482 4870 6534 4922
rect 6546 4870 6598 4922
rect 6610 4870 6662 4922
rect 6674 4870 6726 4922
rect 6738 4870 6790 4922
rect 2412 4768 2464 4820
rect 3884 4632 3936 4684
rect 5448 4632 5500 4684
rect 1584 4607 1636 4616
rect 1584 4573 1593 4607
rect 1593 4573 1627 4607
rect 1627 4573 1636 4607
rect 1584 4564 1636 4573
rect 3148 4564 3200 4616
rect 3792 4564 3844 4616
rect 4068 4564 4120 4616
rect 2504 4496 2556 4548
rect 4068 4428 4120 4480
rect 2658 4326 2710 4378
rect 2722 4326 2774 4378
rect 2786 4326 2838 4378
rect 2850 4326 2902 4378
rect 2914 4326 2966 4378
rect 2978 4326 3030 4378
rect 4158 4326 4210 4378
rect 4222 4326 4274 4378
rect 4286 4326 4338 4378
rect 4350 4326 4402 4378
rect 4414 4326 4466 4378
rect 4478 4326 4530 4378
rect 5658 4326 5710 4378
rect 5722 4326 5774 4378
rect 5786 4326 5838 4378
rect 5850 4326 5902 4378
rect 5914 4326 5966 4378
rect 5978 4326 6030 4378
rect 2412 4224 2464 4276
rect 3240 4224 3292 4276
rect 3332 4156 3384 4208
rect 2504 4088 2556 4140
rect 3240 4088 3292 4140
rect 4528 4088 4580 4140
rect 3240 3884 3292 3936
rect 3792 3884 3844 3936
rect 1918 3782 1970 3834
rect 1982 3782 2034 3834
rect 2046 3782 2098 3834
rect 2110 3782 2162 3834
rect 2174 3782 2226 3834
rect 2238 3782 2290 3834
rect 3418 3782 3470 3834
rect 3482 3782 3534 3834
rect 3546 3782 3598 3834
rect 3610 3782 3662 3834
rect 3674 3782 3726 3834
rect 3738 3782 3790 3834
rect 4918 3782 4970 3834
rect 4982 3782 5034 3834
rect 5046 3782 5098 3834
rect 5110 3782 5162 3834
rect 5174 3782 5226 3834
rect 5238 3782 5290 3834
rect 6418 3782 6470 3834
rect 6482 3782 6534 3834
rect 6546 3782 6598 3834
rect 6610 3782 6662 3834
rect 6674 3782 6726 3834
rect 6738 3782 6790 3834
rect 3884 3723 3936 3732
rect 3884 3689 3893 3723
rect 3893 3689 3927 3723
rect 3927 3689 3936 3723
rect 3884 3680 3936 3689
rect 3056 3612 3108 3664
rect 3148 3544 3200 3596
rect 3884 3544 3936 3596
rect 6184 3544 6236 3596
rect 1584 3519 1636 3528
rect 1584 3485 1593 3519
rect 1593 3485 1627 3519
rect 1627 3485 1636 3519
rect 1584 3476 1636 3485
rect 3332 3476 3384 3528
rect 3240 3408 3292 3460
rect 3976 3340 4028 3392
rect 2658 3238 2710 3290
rect 2722 3238 2774 3290
rect 2786 3238 2838 3290
rect 2850 3238 2902 3290
rect 2914 3238 2966 3290
rect 2978 3238 3030 3290
rect 4158 3238 4210 3290
rect 4222 3238 4274 3290
rect 4286 3238 4338 3290
rect 4350 3238 4402 3290
rect 4414 3238 4466 3290
rect 4478 3238 4530 3290
rect 5658 3238 5710 3290
rect 5722 3238 5774 3290
rect 5786 3238 5838 3290
rect 5850 3238 5902 3290
rect 5914 3238 5966 3290
rect 5978 3238 6030 3290
rect 3976 3136 4028 3188
rect 848 2864 900 2916
rect 3148 3000 3200 3052
rect 4620 3000 4672 3052
rect 1676 2839 1728 2848
rect 1676 2805 1685 2839
rect 1685 2805 1719 2839
rect 1719 2805 1728 2839
rect 1676 2796 1728 2805
rect 4068 2796 4120 2848
rect 1918 2694 1970 2746
rect 1982 2694 2034 2746
rect 2046 2694 2098 2746
rect 2110 2694 2162 2746
rect 2174 2694 2226 2746
rect 2238 2694 2290 2746
rect 3418 2694 3470 2746
rect 3482 2694 3534 2746
rect 3546 2694 3598 2746
rect 3610 2694 3662 2746
rect 3674 2694 3726 2746
rect 3738 2694 3790 2746
rect 4918 2694 4970 2746
rect 4982 2694 5034 2746
rect 5046 2694 5098 2746
rect 5110 2694 5162 2746
rect 5174 2694 5226 2746
rect 5238 2694 5290 2746
rect 6418 2694 6470 2746
rect 6482 2694 6534 2746
rect 6546 2694 6598 2746
rect 6610 2694 6662 2746
rect 6674 2694 6726 2746
rect 6738 2694 6790 2746
rect 1584 2592 1636 2644
rect 3884 2592 3936 2644
rect 4712 2592 4764 2644
rect 3976 2388 4028 2440
rect 5540 2431 5592 2440
rect 5540 2397 5549 2431
rect 5549 2397 5583 2431
rect 5583 2397 5592 2431
rect 5540 2388 5592 2397
rect 2658 2150 2710 2202
rect 2722 2150 2774 2202
rect 2786 2150 2838 2202
rect 2850 2150 2902 2202
rect 2914 2150 2966 2202
rect 2978 2150 3030 2202
rect 4158 2150 4210 2202
rect 4222 2150 4274 2202
rect 4286 2150 4338 2202
rect 4350 2150 4402 2202
rect 4414 2150 4466 2202
rect 4478 2150 4530 2202
rect 5658 2150 5710 2202
rect 5722 2150 5774 2202
rect 5786 2150 5838 2202
rect 5850 2150 5902 2202
rect 5914 2150 5966 2202
rect 5978 2150 6030 2202
<< metal2 >>
rect 1950 9602 2006 10271
rect 5998 9602 6054 10271
rect 1950 9574 2084 9602
rect 1950 9471 2006 9574
rect 1398 8800 1454 8809
rect 1398 8735 1454 8744
rect 1412 7546 1440 8735
rect 1400 7540 1452 7546
rect 1400 7482 1452 7488
rect 2056 7410 2084 9574
rect 5998 9574 6132 9602
rect 5998 9471 6054 9574
rect 2656 7644 3032 7653
rect 2712 7642 2736 7644
rect 2792 7642 2816 7644
rect 2872 7642 2896 7644
rect 2952 7642 2976 7644
rect 2712 7590 2722 7642
rect 2966 7590 2976 7642
rect 2712 7588 2736 7590
rect 2792 7588 2816 7590
rect 2872 7588 2896 7590
rect 2952 7588 2976 7590
rect 2656 7579 3032 7588
rect 4156 7644 4532 7653
rect 4212 7642 4236 7644
rect 4292 7642 4316 7644
rect 4372 7642 4396 7644
rect 4452 7642 4476 7644
rect 4212 7590 4222 7642
rect 4466 7590 4476 7642
rect 4212 7588 4236 7590
rect 4292 7588 4316 7590
rect 4372 7588 4396 7590
rect 4452 7588 4476 7590
rect 4156 7579 4532 7588
rect 5656 7644 6032 7653
rect 5712 7642 5736 7644
rect 5792 7642 5816 7644
rect 5872 7642 5896 7644
rect 5952 7642 5976 7644
rect 5712 7590 5722 7642
rect 5966 7590 5976 7642
rect 5712 7588 5736 7590
rect 5792 7588 5816 7590
rect 5872 7588 5896 7590
rect 5952 7588 5976 7590
rect 5656 7579 6032 7588
rect 2044 7404 2096 7410
rect 2044 7346 2096 7352
rect 3148 7336 3200 7342
rect 3148 7278 3200 7284
rect 1676 7200 1728 7206
rect 1676 7142 1728 7148
rect 3056 7200 3108 7206
rect 3056 7142 3108 7148
rect 1688 6905 1716 7142
rect 1916 7100 2292 7109
rect 1972 7098 1996 7100
rect 2052 7098 2076 7100
rect 2132 7098 2156 7100
rect 2212 7098 2236 7100
rect 1972 7046 1982 7098
rect 2226 7046 2236 7098
rect 1972 7044 1996 7046
rect 2052 7044 2076 7046
rect 2132 7044 2156 7046
rect 2212 7044 2236 7046
rect 1916 7035 2292 7044
rect 1674 6896 1730 6905
rect 1674 6831 1730 6840
rect 2656 6556 3032 6565
rect 2712 6554 2736 6556
rect 2792 6554 2816 6556
rect 2872 6554 2896 6556
rect 2952 6554 2976 6556
rect 2712 6502 2722 6554
rect 2966 6502 2976 6554
rect 2712 6500 2736 6502
rect 2792 6500 2816 6502
rect 2872 6500 2896 6502
rect 2952 6500 2976 6502
rect 2656 6491 3032 6500
rect 2872 6248 2924 6254
rect 2872 6190 2924 6196
rect 1916 6012 2292 6021
rect 1972 6010 1996 6012
rect 2052 6010 2076 6012
rect 2132 6010 2156 6012
rect 2212 6010 2236 6012
rect 1972 5958 1982 6010
rect 2226 5958 2236 6010
rect 1972 5956 1996 5958
rect 2052 5956 2076 5958
rect 2132 5956 2156 5958
rect 2212 5956 2236 5958
rect 1916 5947 2292 5956
rect 1584 5704 1636 5710
rect 1584 5646 1636 5652
rect 846 5128 902 5137
rect 846 5063 902 5072
rect 860 5030 888 5063
rect 848 5024 900 5030
rect 848 4966 900 4972
rect 1596 4622 1624 5646
rect 2884 5574 2912 6190
rect 3068 5914 3096 7142
rect 3056 5908 3108 5914
rect 3056 5850 3108 5856
rect 3056 5772 3108 5778
rect 3056 5714 3108 5720
rect 2872 5568 2924 5574
rect 2872 5510 2924 5516
rect 2656 5468 3032 5477
rect 2712 5466 2736 5468
rect 2792 5466 2816 5468
rect 2872 5466 2896 5468
rect 2952 5466 2976 5468
rect 2712 5414 2722 5466
rect 2966 5414 2976 5466
rect 2712 5412 2736 5414
rect 2792 5412 2816 5414
rect 2872 5412 2896 5414
rect 2952 5412 2976 5414
rect 2656 5403 3032 5412
rect 2412 5228 2464 5234
rect 2412 5170 2464 5176
rect 1916 4924 2292 4933
rect 1972 4922 1996 4924
rect 2052 4922 2076 4924
rect 2132 4922 2156 4924
rect 2212 4922 2236 4924
rect 1972 4870 1982 4922
rect 2226 4870 2236 4922
rect 1972 4868 1996 4870
rect 2052 4868 2076 4870
rect 2132 4868 2156 4870
rect 2212 4868 2236 4870
rect 1916 4859 2292 4868
rect 2424 4826 2452 5170
rect 2412 4820 2464 4826
rect 2412 4762 2464 4768
rect 1584 4616 1636 4622
rect 1584 4558 1636 4564
rect 1596 3534 1624 4558
rect 2424 4282 2452 4762
rect 2504 4548 2556 4554
rect 2504 4490 2556 4496
rect 2412 4276 2464 4282
rect 2412 4218 2464 4224
rect 2516 4146 2544 4490
rect 2656 4380 3032 4389
rect 2712 4378 2736 4380
rect 2792 4378 2816 4380
rect 2872 4378 2896 4380
rect 2952 4378 2976 4380
rect 2712 4326 2722 4378
rect 2966 4326 2976 4378
rect 2712 4324 2736 4326
rect 2792 4324 2816 4326
rect 2872 4324 2896 4326
rect 2952 4324 2976 4326
rect 2656 4315 3032 4324
rect 2504 4140 2556 4146
rect 2504 4082 2556 4088
rect 1916 3836 2292 3845
rect 1972 3834 1996 3836
rect 2052 3834 2076 3836
rect 2132 3834 2156 3836
rect 2212 3834 2236 3836
rect 1972 3782 1982 3834
rect 2226 3782 2236 3834
rect 1972 3780 1996 3782
rect 2052 3780 2076 3782
rect 2132 3780 2156 3782
rect 2212 3780 2236 3782
rect 1916 3771 2292 3780
rect 3068 3670 3096 5714
rect 3160 5370 3188 7278
rect 4068 7268 4120 7274
rect 4068 7210 4120 7216
rect 3416 7100 3792 7109
rect 3472 7098 3496 7100
rect 3552 7098 3576 7100
rect 3632 7098 3656 7100
rect 3712 7098 3736 7100
rect 3472 7046 3482 7098
rect 3726 7046 3736 7098
rect 3472 7044 3496 7046
rect 3552 7044 3576 7046
rect 3632 7044 3656 7046
rect 3712 7044 3736 7046
rect 3416 7035 3792 7044
rect 3884 6384 3936 6390
rect 3884 6326 3936 6332
rect 3416 6012 3792 6021
rect 3472 6010 3496 6012
rect 3552 6010 3576 6012
rect 3632 6010 3656 6012
rect 3712 6010 3736 6012
rect 3472 5958 3482 6010
rect 3726 5958 3736 6010
rect 3472 5956 3496 5958
rect 3552 5956 3576 5958
rect 3632 5956 3656 5958
rect 3712 5956 3736 5958
rect 3416 5947 3792 5956
rect 3896 5914 3924 6326
rect 3976 6180 4028 6186
rect 3976 6122 4028 6128
rect 3884 5908 3936 5914
rect 3884 5850 3936 5856
rect 3988 5794 4016 6122
rect 4080 5914 4108 7210
rect 4916 7100 5292 7109
rect 4972 7098 4996 7100
rect 5052 7098 5076 7100
rect 5132 7098 5156 7100
rect 5212 7098 5236 7100
rect 4972 7046 4982 7098
rect 5226 7046 5236 7098
rect 4972 7044 4996 7046
rect 5052 7044 5076 7046
rect 5132 7044 5156 7046
rect 5212 7044 5236 7046
rect 4916 7035 5292 7044
rect 4712 6724 4764 6730
rect 4712 6666 4764 6672
rect 4156 6556 4532 6565
rect 4212 6554 4236 6556
rect 4292 6554 4316 6556
rect 4372 6554 4396 6556
rect 4452 6554 4476 6556
rect 4212 6502 4222 6554
rect 4466 6502 4476 6554
rect 4212 6500 4236 6502
rect 4292 6500 4316 6502
rect 4372 6500 4396 6502
rect 4452 6500 4476 6502
rect 4156 6491 4532 6500
rect 4068 5908 4120 5914
rect 4068 5850 4120 5856
rect 3988 5766 4108 5794
rect 4080 5642 4108 5766
rect 3332 5636 3384 5642
rect 3332 5578 3384 5584
rect 3976 5636 4028 5642
rect 3976 5578 4028 5584
rect 4068 5636 4120 5642
rect 4068 5578 4120 5584
rect 3148 5364 3200 5370
rect 3148 5306 3200 5312
rect 3160 4706 3188 5306
rect 3344 5234 3372 5578
rect 3884 5568 3936 5574
rect 3884 5510 3936 5516
rect 3332 5228 3384 5234
rect 3332 5170 3384 5176
rect 3896 5114 3924 5510
rect 3988 5302 4016 5578
rect 3976 5296 4028 5302
rect 3976 5238 4028 5244
rect 3896 5086 4016 5114
rect 4080 5098 4108 5578
rect 4156 5468 4532 5477
rect 4212 5466 4236 5468
rect 4292 5466 4316 5468
rect 4372 5466 4396 5468
rect 4452 5466 4476 5468
rect 4212 5414 4222 5466
rect 4466 5414 4476 5466
rect 4212 5412 4236 5414
rect 4292 5412 4316 5414
rect 4372 5412 4396 5414
rect 4452 5412 4476 5414
rect 4156 5403 4532 5412
rect 4620 5160 4672 5166
rect 4620 5102 4672 5108
rect 3416 4924 3792 4933
rect 3472 4922 3496 4924
rect 3552 4922 3576 4924
rect 3632 4922 3656 4924
rect 3712 4922 3736 4924
rect 3472 4870 3482 4922
rect 3726 4870 3736 4922
rect 3472 4868 3496 4870
rect 3552 4868 3576 4870
rect 3632 4868 3656 4870
rect 3712 4868 3736 4870
rect 3416 4859 3792 4868
rect 3160 4678 3280 4706
rect 3148 4616 3200 4622
rect 3148 4558 3200 4564
rect 3056 3664 3108 3670
rect 3056 3606 3108 3612
rect 3160 3602 3188 4558
rect 3252 4282 3280 4678
rect 3884 4684 3936 4690
rect 3884 4626 3936 4632
rect 3792 4616 3844 4622
rect 3792 4558 3844 4564
rect 3240 4276 3292 4282
rect 3240 4218 3292 4224
rect 3332 4208 3384 4214
rect 3332 4150 3384 4156
rect 3240 4140 3292 4146
rect 3240 4082 3292 4088
rect 3252 3942 3280 4082
rect 3240 3936 3292 3942
rect 3240 3878 3292 3884
rect 3148 3596 3200 3602
rect 3148 3538 3200 3544
rect 1584 3528 1636 3534
rect 1584 3470 1636 3476
rect 846 2952 902 2961
rect 846 2887 848 2896
rect 900 2887 902 2896
rect 848 2858 900 2864
rect 1596 2650 1624 3470
rect 3252 3466 3280 3878
rect 3344 3534 3372 4150
rect 3804 3942 3832 4558
rect 3792 3936 3844 3942
rect 3792 3878 3844 3884
rect 3416 3836 3792 3845
rect 3472 3834 3496 3836
rect 3552 3834 3576 3836
rect 3632 3834 3656 3836
rect 3712 3834 3736 3836
rect 3472 3782 3482 3834
rect 3726 3782 3736 3834
rect 3472 3780 3496 3782
rect 3552 3780 3576 3782
rect 3632 3780 3656 3782
rect 3712 3780 3736 3782
rect 3416 3771 3792 3780
rect 3896 3738 3924 4626
rect 3884 3732 3936 3738
rect 3884 3674 3936 3680
rect 3988 3618 4016 5086
rect 4068 5092 4120 5098
rect 4068 5034 4120 5040
rect 4080 4622 4108 5034
rect 4068 4616 4120 4622
rect 4068 4558 4120 4564
rect 4068 4480 4120 4486
rect 4068 4422 4120 4428
rect 3896 3602 4016 3618
rect 3884 3596 4016 3602
rect 3936 3590 4016 3596
rect 3884 3538 3936 3544
rect 3332 3528 3384 3534
rect 3332 3470 3384 3476
rect 3240 3460 3292 3466
rect 3240 3402 3292 3408
rect 2656 3292 3032 3301
rect 2712 3290 2736 3292
rect 2792 3290 2816 3292
rect 2872 3290 2896 3292
rect 2952 3290 2976 3292
rect 2712 3238 2722 3290
rect 2966 3238 2976 3290
rect 2712 3236 2736 3238
rect 2792 3236 2816 3238
rect 2872 3236 2896 3238
rect 2952 3236 2976 3238
rect 2656 3227 3032 3236
rect 3252 3074 3280 3402
rect 3160 3058 3280 3074
rect 3148 3052 3280 3058
rect 3200 3046 3280 3052
rect 3148 2994 3200 3000
rect 1676 2848 1728 2854
rect 1676 2790 1728 2796
rect 1584 2644 1636 2650
rect 1584 2586 1636 2592
rect 1688 1193 1716 2790
rect 1916 2748 2292 2757
rect 1972 2746 1996 2748
rect 2052 2746 2076 2748
rect 2132 2746 2156 2748
rect 2212 2746 2236 2748
rect 1972 2694 1982 2746
rect 2226 2694 2236 2746
rect 1972 2692 1996 2694
rect 2052 2692 2076 2694
rect 2132 2692 2156 2694
rect 2212 2692 2236 2694
rect 1916 2683 2292 2692
rect 3416 2748 3792 2757
rect 3472 2746 3496 2748
rect 3552 2746 3576 2748
rect 3632 2746 3656 2748
rect 3712 2746 3736 2748
rect 3472 2694 3482 2746
rect 3726 2694 3736 2746
rect 3472 2692 3496 2694
rect 3552 2692 3576 2694
rect 3632 2692 3656 2694
rect 3712 2692 3736 2694
rect 3416 2683 3792 2692
rect 3896 2650 3924 3538
rect 3976 3392 4028 3398
rect 3976 3334 4028 3340
rect 3988 3194 4016 3334
rect 3976 3188 4028 3194
rect 3976 3130 4028 3136
rect 4080 2854 4108 4422
rect 4156 4380 4532 4389
rect 4212 4378 4236 4380
rect 4292 4378 4316 4380
rect 4372 4378 4396 4380
rect 4452 4378 4476 4380
rect 4212 4326 4222 4378
rect 4466 4326 4476 4378
rect 4212 4324 4236 4326
rect 4292 4324 4316 4326
rect 4372 4324 4396 4326
rect 4452 4324 4476 4326
rect 4156 4315 4532 4324
rect 4528 4140 4580 4146
rect 4528 4082 4580 4088
rect 4540 4026 4568 4082
rect 4632 4026 4660 5102
rect 4540 3998 4660 4026
rect 4156 3292 4532 3301
rect 4212 3290 4236 3292
rect 4292 3290 4316 3292
rect 4372 3290 4396 3292
rect 4452 3290 4476 3292
rect 4212 3238 4222 3290
rect 4466 3238 4476 3290
rect 4212 3236 4236 3238
rect 4292 3236 4316 3238
rect 4372 3236 4396 3238
rect 4452 3236 4476 3238
rect 4156 3227 4532 3236
rect 4632 3058 4660 3998
rect 4620 3052 4672 3058
rect 4620 2994 4672 3000
rect 4068 2848 4120 2854
rect 4068 2790 4120 2796
rect 4724 2650 4752 6666
rect 5656 6556 6032 6565
rect 5712 6554 5736 6556
rect 5792 6554 5816 6556
rect 5872 6554 5896 6556
rect 5952 6554 5976 6556
rect 5712 6502 5722 6554
rect 5966 6502 5976 6554
rect 5712 6500 5736 6502
rect 5792 6500 5816 6502
rect 5872 6500 5896 6502
rect 5952 6500 5976 6502
rect 5656 6491 6032 6500
rect 5448 6112 5500 6118
rect 5448 6054 5500 6060
rect 4916 6012 5292 6021
rect 4972 6010 4996 6012
rect 5052 6010 5076 6012
rect 5132 6010 5156 6012
rect 5212 6010 5236 6012
rect 4972 5958 4982 6010
rect 5226 5958 5236 6010
rect 4972 5956 4996 5958
rect 5052 5956 5076 5958
rect 5132 5956 5156 5958
rect 5212 5956 5236 5958
rect 4916 5947 5292 5956
rect 5460 5234 5488 6054
rect 6104 5681 6132 9574
rect 6416 7100 6792 7109
rect 6472 7098 6496 7100
rect 6552 7098 6576 7100
rect 6632 7098 6656 7100
rect 6712 7098 6736 7100
rect 6472 7046 6482 7098
rect 6726 7046 6736 7098
rect 6472 7044 6496 7046
rect 6552 7044 6576 7046
rect 6632 7044 6656 7046
rect 6712 7044 6736 7046
rect 6416 7035 6792 7044
rect 6184 6656 6236 6662
rect 6184 6598 6236 6604
rect 6196 5778 6224 6598
rect 6416 6012 6792 6021
rect 6472 6010 6496 6012
rect 6552 6010 6576 6012
rect 6632 6010 6656 6012
rect 6712 6010 6736 6012
rect 6472 5958 6482 6010
rect 6726 5958 6736 6010
rect 6472 5956 6496 5958
rect 6552 5956 6576 5958
rect 6632 5956 6656 5958
rect 6712 5956 6736 5958
rect 6416 5947 6792 5956
rect 6184 5772 6236 5778
rect 6184 5714 6236 5720
rect 6090 5672 6146 5681
rect 6090 5607 6146 5616
rect 5656 5468 6032 5477
rect 5712 5466 5736 5468
rect 5792 5466 5816 5468
rect 5872 5466 5896 5468
rect 5952 5466 5976 5468
rect 5712 5414 5722 5466
rect 5966 5414 5976 5466
rect 5712 5412 5736 5414
rect 5792 5412 5816 5414
rect 5872 5412 5896 5414
rect 5952 5412 5976 5414
rect 5656 5403 6032 5412
rect 5448 5228 5500 5234
rect 5448 5170 5500 5176
rect 5448 5092 5500 5098
rect 5448 5034 5500 5040
rect 4916 4924 5292 4933
rect 4972 4922 4996 4924
rect 5052 4922 5076 4924
rect 5132 4922 5156 4924
rect 5212 4922 5236 4924
rect 4972 4870 4982 4922
rect 5226 4870 5236 4922
rect 4972 4868 4996 4870
rect 5052 4868 5076 4870
rect 5132 4868 5156 4870
rect 5212 4868 5236 4870
rect 4916 4859 5292 4868
rect 5460 4690 5488 5034
rect 5448 4684 5500 4690
rect 5448 4626 5500 4632
rect 5656 4380 6032 4389
rect 5712 4378 5736 4380
rect 5792 4378 5816 4380
rect 5872 4378 5896 4380
rect 5952 4378 5976 4380
rect 5712 4326 5722 4378
rect 5966 4326 5976 4378
rect 5712 4324 5736 4326
rect 5792 4324 5816 4326
rect 5872 4324 5896 4326
rect 5952 4324 5976 4326
rect 5656 4315 6032 4324
rect 4916 3836 5292 3845
rect 4972 3834 4996 3836
rect 5052 3834 5076 3836
rect 5132 3834 5156 3836
rect 5212 3834 5236 3836
rect 4972 3782 4982 3834
rect 5226 3782 5236 3834
rect 4972 3780 4996 3782
rect 5052 3780 5076 3782
rect 5132 3780 5156 3782
rect 5212 3780 5236 3782
rect 4916 3771 5292 3780
rect 6196 3602 6224 5714
rect 6920 5228 6972 5234
rect 6920 5170 6972 5176
rect 6932 5001 6960 5170
rect 6918 4992 6974 5001
rect 6416 4924 6792 4933
rect 6918 4927 6974 4936
rect 6472 4922 6496 4924
rect 6552 4922 6576 4924
rect 6632 4922 6656 4924
rect 6712 4922 6736 4924
rect 6472 4870 6482 4922
rect 6726 4870 6736 4922
rect 6472 4868 6496 4870
rect 6552 4868 6576 4870
rect 6632 4868 6656 4870
rect 6712 4868 6736 4870
rect 6416 4859 6792 4868
rect 6416 3836 6792 3845
rect 6472 3834 6496 3836
rect 6552 3834 6576 3836
rect 6632 3834 6656 3836
rect 6712 3834 6736 3836
rect 6472 3782 6482 3834
rect 6726 3782 6736 3834
rect 6472 3780 6496 3782
rect 6552 3780 6576 3782
rect 6632 3780 6656 3782
rect 6712 3780 6736 3782
rect 6416 3771 6792 3780
rect 6184 3596 6236 3602
rect 6184 3538 6236 3544
rect 5656 3292 6032 3301
rect 5712 3290 5736 3292
rect 5792 3290 5816 3292
rect 5872 3290 5896 3292
rect 5952 3290 5976 3292
rect 5712 3238 5722 3290
rect 5966 3238 5976 3290
rect 5712 3236 5736 3238
rect 5792 3236 5816 3238
rect 5872 3236 5896 3238
rect 5952 3236 5976 3238
rect 5656 3227 6032 3236
rect 4916 2748 5292 2757
rect 4972 2746 4996 2748
rect 5052 2746 5076 2748
rect 5132 2746 5156 2748
rect 5212 2746 5236 2748
rect 4972 2694 4982 2746
rect 5226 2694 5236 2746
rect 4972 2692 4996 2694
rect 5052 2692 5076 2694
rect 5132 2692 5156 2694
rect 5212 2692 5236 2694
rect 4916 2683 5292 2692
rect 6416 2748 6792 2757
rect 6472 2746 6496 2748
rect 6552 2746 6576 2748
rect 6632 2746 6656 2748
rect 6712 2746 6736 2748
rect 6472 2694 6482 2746
rect 6726 2694 6736 2746
rect 6472 2692 6496 2694
rect 6552 2692 6576 2694
rect 6632 2692 6656 2694
rect 6712 2692 6736 2694
rect 5538 2680 5594 2689
rect 6416 2683 6792 2692
rect 3884 2644 3936 2650
rect 3884 2586 3936 2592
rect 4712 2644 4764 2650
rect 5538 2615 5594 2624
rect 4712 2586 4764 2592
rect 5552 2446 5580 2615
rect 3976 2440 4028 2446
rect 3976 2382 4028 2388
rect 5540 2440 5592 2446
rect 5540 2382 5592 2388
rect 2656 2204 3032 2213
rect 2712 2202 2736 2204
rect 2792 2202 2816 2204
rect 2872 2202 2896 2204
rect 2952 2202 2976 2204
rect 2712 2150 2722 2202
rect 2966 2150 2976 2202
rect 2712 2148 2736 2150
rect 2792 2148 2816 2150
rect 2872 2148 2896 2150
rect 2952 2148 2976 2150
rect 2656 2139 3032 2148
rect 1674 1184 1730 1193
rect 1674 1119 1730 1128
rect 3988 800 4016 2382
rect 4156 2204 4532 2213
rect 4212 2202 4236 2204
rect 4292 2202 4316 2204
rect 4372 2202 4396 2204
rect 4452 2202 4476 2204
rect 4212 2150 4222 2202
rect 4466 2150 4476 2202
rect 4212 2148 4236 2150
rect 4292 2148 4316 2150
rect 4372 2148 4396 2150
rect 4452 2148 4476 2150
rect 4156 2139 4532 2148
rect 5656 2204 6032 2213
rect 5712 2202 5736 2204
rect 5792 2202 5816 2204
rect 5872 2202 5896 2204
rect 5952 2202 5976 2204
rect 5712 2150 5722 2202
rect 5966 2150 5976 2202
rect 5712 2148 5736 2150
rect 5792 2148 5816 2150
rect 5872 2148 5896 2150
rect 5952 2148 5976 2150
rect 5656 2139 6032 2148
rect 3974 0 4030 800
<< via2 >>
rect 1398 8744 1454 8800
rect 2656 7642 2712 7644
rect 2736 7642 2792 7644
rect 2816 7642 2872 7644
rect 2896 7642 2952 7644
rect 2976 7642 3032 7644
rect 2656 7590 2658 7642
rect 2658 7590 2710 7642
rect 2710 7590 2712 7642
rect 2736 7590 2774 7642
rect 2774 7590 2786 7642
rect 2786 7590 2792 7642
rect 2816 7590 2838 7642
rect 2838 7590 2850 7642
rect 2850 7590 2872 7642
rect 2896 7590 2902 7642
rect 2902 7590 2914 7642
rect 2914 7590 2952 7642
rect 2976 7590 2978 7642
rect 2978 7590 3030 7642
rect 3030 7590 3032 7642
rect 2656 7588 2712 7590
rect 2736 7588 2792 7590
rect 2816 7588 2872 7590
rect 2896 7588 2952 7590
rect 2976 7588 3032 7590
rect 4156 7642 4212 7644
rect 4236 7642 4292 7644
rect 4316 7642 4372 7644
rect 4396 7642 4452 7644
rect 4476 7642 4532 7644
rect 4156 7590 4158 7642
rect 4158 7590 4210 7642
rect 4210 7590 4212 7642
rect 4236 7590 4274 7642
rect 4274 7590 4286 7642
rect 4286 7590 4292 7642
rect 4316 7590 4338 7642
rect 4338 7590 4350 7642
rect 4350 7590 4372 7642
rect 4396 7590 4402 7642
rect 4402 7590 4414 7642
rect 4414 7590 4452 7642
rect 4476 7590 4478 7642
rect 4478 7590 4530 7642
rect 4530 7590 4532 7642
rect 4156 7588 4212 7590
rect 4236 7588 4292 7590
rect 4316 7588 4372 7590
rect 4396 7588 4452 7590
rect 4476 7588 4532 7590
rect 5656 7642 5712 7644
rect 5736 7642 5792 7644
rect 5816 7642 5872 7644
rect 5896 7642 5952 7644
rect 5976 7642 6032 7644
rect 5656 7590 5658 7642
rect 5658 7590 5710 7642
rect 5710 7590 5712 7642
rect 5736 7590 5774 7642
rect 5774 7590 5786 7642
rect 5786 7590 5792 7642
rect 5816 7590 5838 7642
rect 5838 7590 5850 7642
rect 5850 7590 5872 7642
rect 5896 7590 5902 7642
rect 5902 7590 5914 7642
rect 5914 7590 5952 7642
rect 5976 7590 5978 7642
rect 5978 7590 6030 7642
rect 6030 7590 6032 7642
rect 5656 7588 5712 7590
rect 5736 7588 5792 7590
rect 5816 7588 5872 7590
rect 5896 7588 5952 7590
rect 5976 7588 6032 7590
rect 1916 7098 1972 7100
rect 1996 7098 2052 7100
rect 2076 7098 2132 7100
rect 2156 7098 2212 7100
rect 2236 7098 2292 7100
rect 1916 7046 1918 7098
rect 1918 7046 1970 7098
rect 1970 7046 1972 7098
rect 1996 7046 2034 7098
rect 2034 7046 2046 7098
rect 2046 7046 2052 7098
rect 2076 7046 2098 7098
rect 2098 7046 2110 7098
rect 2110 7046 2132 7098
rect 2156 7046 2162 7098
rect 2162 7046 2174 7098
rect 2174 7046 2212 7098
rect 2236 7046 2238 7098
rect 2238 7046 2290 7098
rect 2290 7046 2292 7098
rect 1916 7044 1972 7046
rect 1996 7044 2052 7046
rect 2076 7044 2132 7046
rect 2156 7044 2212 7046
rect 2236 7044 2292 7046
rect 1674 6840 1730 6896
rect 2656 6554 2712 6556
rect 2736 6554 2792 6556
rect 2816 6554 2872 6556
rect 2896 6554 2952 6556
rect 2976 6554 3032 6556
rect 2656 6502 2658 6554
rect 2658 6502 2710 6554
rect 2710 6502 2712 6554
rect 2736 6502 2774 6554
rect 2774 6502 2786 6554
rect 2786 6502 2792 6554
rect 2816 6502 2838 6554
rect 2838 6502 2850 6554
rect 2850 6502 2872 6554
rect 2896 6502 2902 6554
rect 2902 6502 2914 6554
rect 2914 6502 2952 6554
rect 2976 6502 2978 6554
rect 2978 6502 3030 6554
rect 3030 6502 3032 6554
rect 2656 6500 2712 6502
rect 2736 6500 2792 6502
rect 2816 6500 2872 6502
rect 2896 6500 2952 6502
rect 2976 6500 3032 6502
rect 1916 6010 1972 6012
rect 1996 6010 2052 6012
rect 2076 6010 2132 6012
rect 2156 6010 2212 6012
rect 2236 6010 2292 6012
rect 1916 5958 1918 6010
rect 1918 5958 1970 6010
rect 1970 5958 1972 6010
rect 1996 5958 2034 6010
rect 2034 5958 2046 6010
rect 2046 5958 2052 6010
rect 2076 5958 2098 6010
rect 2098 5958 2110 6010
rect 2110 5958 2132 6010
rect 2156 5958 2162 6010
rect 2162 5958 2174 6010
rect 2174 5958 2212 6010
rect 2236 5958 2238 6010
rect 2238 5958 2290 6010
rect 2290 5958 2292 6010
rect 1916 5956 1972 5958
rect 1996 5956 2052 5958
rect 2076 5956 2132 5958
rect 2156 5956 2212 5958
rect 2236 5956 2292 5958
rect 846 5072 902 5128
rect 2656 5466 2712 5468
rect 2736 5466 2792 5468
rect 2816 5466 2872 5468
rect 2896 5466 2952 5468
rect 2976 5466 3032 5468
rect 2656 5414 2658 5466
rect 2658 5414 2710 5466
rect 2710 5414 2712 5466
rect 2736 5414 2774 5466
rect 2774 5414 2786 5466
rect 2786 5414 2792 5466
rect 2816 5414 2838 5466
rect 2838 5414 2850 5466
rect 2850 5414 2872 5466
rect 2896 5414 2902 5466
rect 2902 5414 2914 5466
rect 2914 5414 2952 5466
rect 2976 5414 2978 5466
rect 2978 5414 3030 5466
rect 3030 5414 3032 5466
rect 2656 5412 2712 5414
rect 2736 5412 2792 5414
rect 2816 5412 2872 5414
rect 2896 5412 2952 5414
rect 2976 5412 3032 5414
rect 1916 4922 1972 4924
rect 1996 4922 2052 4924
rect 2076 4922 2132 4924
rect 2156 4922 2212 4924
rect 2236 4922 2292 4924
rect 1916 4870 1918 4922
rect 1918 4870 1970 4922
rect 1970 4870 1972 4922
rect 1996 4870 2034 4922
rect 2034 4870 2046 4922
rect 2046 4870 2052 4922
rect 2076 4870 2098 4922
rect 2098 4870 2110 4922
rect 2110 4870 2132 4922
rect 2156 4870 2162 4922
rect 2162 4870 2174 4922
rect 2174 4870 2212 4922
rect 2236 4870 2238 4922
rect 2238 4870 2290 4922
rect 2290 4870 2292 4922
rect 1916 4868 1972 4870
rect 1996 4868 2052 4870
rect 2076 4868 2132 4870
rect 2156 4868 2212 4870
rect 2236 4868 2292 4870
rect 2656 4378 2712 4380
rect 2736 4378 2792 4380
rect 2816 4378 2872 4380
rect 2896 4378 2952 4380
rect 2976 4378 3032 4380
rect 2656 4326 2658 4378
rect 2658 4326 2710 4378
rect 2710 4326 2712 4378
rect 2736 4326 2774 4378
rect 2774 4326 2786 4378
rect 2786 4326 2792 4378
rect 2816 4326 2838 4378
rect 2838 4326 2850 4378
rect 2850 4326 2872 4378
rect 2896 4326 2902 4378
rect 2902 4326 2914 4378
rect 2914 4326 2952 4378
rect 2976 4326 2978 4378
rect 2978 4326 3030 4378
rect 3030 4326 3032 4378
rect 2656 4324 2712 4326
rect 2736 4324 2792 4326
rect 2816 4324 2872 4326
rect 2896 4324 2952 4326
rect 2976 4324 3032 4326
rect 1916 3834 1972 3836
rect 1996 3834 2052 3836
rect 2076 3834 2132 3836
rect 2156 3834 2212 3836
rect 2236 3834 2292 3836
rect 1916 3782 1918 3834
rect 1918 3782 1970 3834
rect 1970 3782 1972 3834
rect 1996 3782 2034 3834
rect 2034 3782 2046 3834
rect 2046 3782 2052 3834
rect 2076 3782 2098 3834
rect 2098 3782 2110 3834
rect 2110 3782 2132 3834
rect 2156 3782 2162 3834
rect 2162 3782 2174 3834
rect 2174 3782 2212 3834
rect 2236 3782 2238 3834
rect 2238 3782 2290 3834
rect 2290 3782 2292 3834
rect 1916 3780 1972 3782
rect 1996 3780 2052 3782
rect 2076 3780 2132 3782
rect 2156 3780 2212 3782
rect 2236 3780 2292 3782
rect 3416 7098 3472 7100
rect 3496 7098 3552 7100
rect 3576 7098 3632 7100
rect 3656 7098 3712 7100
rect 3736 7098 3792 7100
rect 3416 7046 3418 7098
rect 3418 7046 3470 7098
rect 3470 7046 3472 7098
rect 3496 7046 3534 7098
rect 3534 7046 3546 7098
rect 3546 7046 3552 7098
rect 3576 7046 3598 7098
rect 3598 7046 3610 7098
rect 3610 7046 3632 7098
rect 3656 7046 3662 7098
rect 3662 7046 3674 7098
rect 3674 7046 3712 7098
rect 3736 7046 3738 7098
rect 3738 7046 3790 7098
rect 3790 7046 3792 7098
rect 3416 7044 3472 7046
rect 3496 7044 3552 7046
rect 3576 7044 3632 7046
rect 3656 7044 3712 7046
rect 3736 7044 3792 7046
rect 3416 6010 3472 6012
rect 3496 6010 3552 6012
rect 3576 6010 3632 6012
rect 3656 6010 3712 6012
rect 3736 6010 3792 6012
rect 3416 5958 3418 6010
rect 3418 5958 3470 6010
rect 3470 5958 3472 6010
rect 3496 5958 3534 6010
rect 3534 5958 3546 6010
rect 3546 5958 3552 6010
rect 3576 5958 3598 6010
rect 3598 5958 3610 6010
rect 3610 5958 3632 6010
rect 3656 5958 3662 6010
rect 3662 5958 3674 6010
rect 3674 5958 3712 6010
rect 3736 5958 3738 6010
rect 3738 5958 3790 6010
rect 3790 5958 3792 6010
rect 3416 5956 3472 5958
rect 3496 5956 3552 5958
rect 3576 5956 3632 5958
rect 3656 5956 3712 5958
rect 3736 5956 3792 5958
rect 4916 7098 4972 7100
rect 4996 7098 5052 7100
rect 5076 7098 5132 7100
rect 5156 7098 5212 7100
rect 5236 7098 5292 7100
rect 4916 7046 4918 7098
rect 4918 7046 4970 7098
rect 4970 7046 4972 7098
rect 4996 7046 5034 7098
rect 5034 7046 5046 7098
rect 5046 7046 5052 7098
rect 5076 7046 5098 7098
rect 5098 7046 5110 7098
rect 5110 7046 5132 7098
rect 5156 7046 5162 7098
rect 5162 7046 5174 7098
rect 5174 7046 5212 7098
rect 5236 7046 5238 7098
rect 5238 7046 5290 7098
rect 5290 7046 5292 7098
rect 4916 7044 4972 7046
rect 4996 7044 5052 7046
rect 5076 7044 5132 7046
rect 5156 7044 5212 7046
rect 5236 7044 5292 7046
rect 4156 6554 4212 6556
rect 4236 6554 4292 6556
rect 4316 6554 4372 6556
rect 4396 6554 4452 6556
rect 4476 6554 4532 6556
rect 4156 6502 4158 6554
rect 4158 6502 4210 6554
rect 4210 6502 4212 6554
rect 4236 6502 4274 6554
rect 4274 6502 4286 6554
rect 4286 6502 4292 6554
rect 4316 6502 4338 6554
rect 4338 6502 4350 6554
rect 4350 6502 4372 6554
rect 4396 6502 4402 6554
rect 4402 6502 4414 6554
rect 4414 6502 4452 6554
rect 4476 6502 4478 6554
rect 4478 6502 4530 6554
rect 4530 6502 4532 6554
rect 4156 6500 4212 6502
rect 4236 6500 4292 6502
rect 4316 6500 4372 6502
rect 4396 6500 4452 6502
rect 4476 6500 4532 6502
rect 4156 5466 4212 5468
rect 4236 5466 4292 5468
rect 4316 5466 4372 5468
rect 4396 5466 4452 5468
rect 4476 5466 4532 5468
rect 4156 5414 4158 5466
rect 4158 5414 4210 5466
rect 4210 5414 4212 5466
rect 4236 5414 4274 5466
rect 4274 5414 4286 5466
rect 4286 5414 4292 5466
rect 4316 5414 4338 5466
rect 4338 5414 4350 5466
rect 4350 5414 4372 5466
rect 4396 5414 4402 5466
rect 4402 5414 4414 5466
rect 4414 5414 4452 5466
rect 4476 5414 4478 5466
rect 4478 5414 4530 5466
rect 4530 5414 4532 5466
rect 4156 5412 4212 5414
rect 4236 5412 4292 5414
rect 4316 5412 4372 5414
rect 4396 5412 4452 5414
rect 4476 5412 4532 5414
rect 3416 4922 3472 4924
rect 3496 4922 3552 4924
rect 3576 4922 3632 4924
rect 3656 4922 3712 4924
rect 3736 4922 3792 4924
rect 3416 4870 3418 4922
rect 3418 4870 3470 4922
rect 3470 4870 3472 4922
rect 3496 4870 3534 4922
rect 3534 4870 3546 4922
rect 3546 4870 3552 4922
rect 3576 4870 3598 4922
rect 3598 4870 3610 4922
rect 3610 4870 3632 4922
rect 3656 4870 3662 4922
rect 3662 4870 3674 4922
rect 3674 4870 3712 4922
rect 3736 4870 3738 4922
rect 3738 4870 3790 4922
rect 3790 4870 3792 4922
rect 3416 4868 3472 4870
rect 3496 4868 3552 4870
rect 3576 4868 3632 4870
rect 3656 4868 3712 4870
rect 3736 4868 3792 4870
rect 846 2916 902 2952
rect 846 2896 848 2916
rect 848 2896 900 2916
rect 900 2896 902 2916
rect 3416 3834 3472 3836
rect 3496 3834 3552 3836
rect 3576 3834 3632 3836
rect 3656 3834 3712 3836
rect 3736 3834 3792 3836
rect 3416 3782 3418 3834
rect 3418 3782 3470 3834
rect 3470 3782 3472 3834
rect 3496 3782 3534 3834
rect 3534 3782 3546 3834
rect 3546 3782 3552 3834
rect 3576 3782 3598 3834
rect 3598 3782 3610 3834
rect 3610 3782 3632 3834
rect 3656 3782 3662 3834
rect 3662 3782 3674 3834
rect 3674 3782 3712 3834
rect 3736 3782 3738 3834
rect 3738 3782 3790 3834
rect 3790 3782 3792 3834
rect 3416 3780 3472 3782
rect 3496 3780 3552 3782
rect 3576 3780 3632 3782
rect 3656 3780 3712 3782
rect 3736 3780 3792 3782
rect 2656 3290 2712 3292
rect 2736 3290 2792 3292
rect 2816 3290 2872 3292
rect 2896 3290 2952 3292
rect 2976 3290 3032 3292
rect 2656 3238 2658 3290
rect 2658 3238 2710 3290
rect 2710 3238 2712 3290
rect 2736 3238 2774 3290
rect 2774 3238 2786 3290
rect 2786 3238 2792 3290
rect 2816 3238 2838 3290
rect 2838 3238 2850 3290
rect 2850 3238 2872 3290
rect 2896 3238 2902 3290
rect 2902 3238 2914 3290
rect 2914 3238 2952 3290
rect 2976 3238 2978 3290
rect 2978 3238 3030 3290
rect 3030 3238 3032 3290
rect 2656 3236 2712 3238
rect 2736 3236 2792 3238
rect 2816 3236 2872 3238
rect 2896 3236 2952 3238
rect 2976 3236 3032 3238
rect 1916 2746 1972 2748
rect 1996 2746 2052 2748
rect 2076 2746 2132 2748
rect 2156 2746 2212 2748
rect 2236 2746 2292 2748
rect 1916 2694 1918 2746
rect 1918 2694 1970 2746
rect 1970 2694 1972 2746
rect 1996 2694 2034 2746
rect 2034 2694 2046 2746
rect 2046 2694 2052 2746
rect 2076 2694 2098 2746
rect 2098 2694 2110 2746
rect 2110 2694 2132 2746
rect 2156 2694 2162 2746
rect 2162 2694 2174 2746
rect 2174 2694 2212 2746
rect 2236 2694 2238 2746
rect 2238 2694 2290 2746
rect 2290 2694 2292 2746
rect 1916 2692 1972 2694
rect 1996 2692 2052 2694
rect 2076 2692 2132 2694
rect 2156 2692 2212 2694
rect 2236 2692 2292 2694
rect 3416 2746 3472 2748
rect 3496 2746 3552 2748
rect 3576 2746 3632 2748
rect 3656 2746 3712 2748
rect 3736 2746 3792 2748
rect 3416 2694 3418 2746
rect 3418 2694 3470 2746
rect 3470 2694 3472 2746
rect 3496 2694 3534 2746
rect 3534 2694 3546 2746
rect 3546 2694 3552 2746
rect 3576 2694 3598 2746
rect 3598 2694 3610 2746
rect 3610 2694 3632 2746
rect 3656 2694 3662 2746
rect 3662 2694 3674 2746
rect 3674 2694 3712 2746
rect 3736 2694 3738 2746
rect 3738 2694 3790 2746
rect 3790 2694 3792 2746
rect 3416 2692 3472 2694
rect 3496 2692 3552 2694
rect 3576 2692 3632 2694
rect 3656 2692 3712 2694
rect 3736 2692 3792 2694
rect 4156 4378 4212 4380
rect 4236 4378 4292 4380
rect 4316 4378 4372 4380
rect 4396 4378 4452 4380
rect 4476 4378 4532 4380
rect 4156 4326 4158 4378
rect 4158 4326 4210 4378
rect 4210 4326 4212 4378
rect 4236 4326 4274 4378
rect 4274 4326 4286 4378
rect 4286 4326 4292 4378
rect 4316 4326 4338 4378
rect 4338 4326 4350 4378
rect 4350 4326 4372 4378
rect 4396 4326 4402 4378
rect 4402 4326 4414 4378
rect 4414 4326 4452 4378
rect 4476 4326 4478 4378
rect 4478 4326 4530 4378
rect 4530 4326 4532 4378
rect 4156 4324 4212 4326
rect 4236 4324 4292 4326
rect 4316 4324 4372 4326
rect 4396 4324 4452 4326
rect 4476 4324 4532 4326
rect 4156 3290 4212 3292
rect 4236 3290 4292 3292
rect 4316 3290 4372 3292
rect 4396 3290 4452 3292
rect 4476 3290 4532 3292
rect 4156 3238 4158 3290
rect 4158 3238 4210 3290
rect 4210 3238 4212 3290
rect 4236 3238 4274 3290
rect 4274 3238 4286 3290
rect 4286 3238 4292 3290
rect 4316 3238 4338 3290
rect 4338 3238 4350 3290
rect 4350 3238 4372 3290
rect 4396 3238 4402 3290
rect 4402 3238 4414 3290
rect 4414 3238 4452 3290
rect 4476 3238 4478 3290
rect 4478 3238 4530 3290
rect 4530 3238 4532 3290
rect 4156 3236 4212 3238
rect 4236 3236 4292 3238
rect 4316 3236 4372 3238
rect 4396 3236 4452 3238
rect 4476 3236 4532 3238
rect 5656 6554 5712 6556
rect 5736 6554 5792 6556
rect 5816 6554 5872 6556
rect 5896 6554 5952 6556
rect 5976 6554 6032 6556
rect 5656 6502 5658 6554
rect 5658 6502 5710 6554
rect 5710 6502 5712 6554
rect 5736 6502 5774 6554
rect 5774 6502 5786 6554
rect 5786 6502 5792 6554
rect 5816 6502 5838 6554
rect 5838 6502 5850 6554
rect 5850 6502 5872 6554
rect 5896 6502 5902 6554
rect 5902 6502 5914 6554
rect 5914 6502 5952 6554
rect 5976 6502 5978 6554
rect 5978 6502 6030 6554
rect 6030 6502 6032 6554
rect 5656 6500 5712 6502
rect 5736 6500 5792 6502
rect 5816 6500 5872 6502
rect 5896 6500 5952 6502
rect 5976 6500 6032 6502
rect 4916 6010 4972 6012
rect 4996 6010 5052 6012
rect 5076 6010 5132 6012
rect 5156 6010 5212 6012
rect 5236 6010 5292 6012
rect 4916 5958 4918 6010
rect 4918 5958 4970 6010
rect 4970 5958 4972 6010
rect 4996 5958 5034 6010
rect 5034 5958 5046 6010
rect 5046 5958 5052 6010
rect 5076 5958 5098 6010
rect 5098 5958 5110 6010
rect 5110 5958 5132 6010
rect 5156 5958 5162 6010
rect 5162 5958 5174 6010
rect 5174 5958 5212 6010
rect 5236 5958 5238 6010
rect 5238 5958 5290 6010
rect 5290 5958 5292 6010
rect 4916 5956 4972 5958
rect 4996 5956 5052 5958
rect 5076 5956 5132 5958
rect 5156 5956 5212 5958
rect 5236 5956 5292 5958
rect 6416 7098 6472 7100
rect 6496 7098 6552 7100
rect 6576 7098 6632 7100
rect 6656 7098 6712 7100
rect 6736 7098 6792 7100
rect 6416 7046 6418 7098
rect 6418 7046 6470 7098
rect 6470 7046 6472 7098
rect 6496 7046 6534 7098
rect 6534 7046 6546 7098
rect 6546 7046 6552 7098
rect 6576 7046 6598 7098
rect 6598 7046 6610 7098
rect 6610 7046 6632 7098
rect 6656 7046 6662 7098
rect 6662 7046 6674 7098
rect 6674 7046 6712 7098
rect 6736 7046 6738 7098
rect 6738 7046 6790 7098
rect 6790 7046 6792 7098
rect 6416 7044 6472 7046
rect 6496 7044 6552 7046
rect 6576 7044 6632 7046
rect 6656 7044 6712 7046
rect 6736 7044 6792 7046
rect 6416 6010 6472 6012
rect 6496 6010 6552 6012
rect 6576 6010 6632 6012
rect 6656 6010 6712 6012
rect 6736 6010 6792 6012
rect 6416 5958 6418 6010
rect 6418 5958 6470 6010
rect 6470 5958 6472 6010
rect 6496 5958 6534 6010
rect 6534 5958 6546 6010
rect 6546 5958 6552 6010
rect 6576 5958 6598 6010
rect 6598 5958 6610 6010
rect 6610 5958 6632 6010
rect 6656 5958 6662 6010
rect 6662 5958 6674 6010
rect 6674 5958 6712 6010
rect 6736 5958 6738 6010
rect 6738 5958 6790 6010
rect 6790 5958 6792 6010
rect 6416 5956 6472 5958
rect 6496 5956 6552 5958
rect 6576 5956 6632 5958
rect 6656 5956 6712 5958
rect 6736 5956 6792 5958
rect 6090 5616 6146 5672
rect 5656 5466 5712 5468
rect 5736 5466 5792 5468
rect 5816 5466 5872 5468
rect 5896 5466 5952 5468
rect 5976 5466 6032 5468
rect 5656 5414 5658 5466
rect 5658 5414 5710 5466
rect 5710 5414 5712 5466
rect 5736 5414 5774 5466
rect 5774 5414 5786 5466
rect 5786 5414 5792 5466
rect 5816 5414 5838 5466
rect 5838 5414 5850 5466
rect 5850 5414 5872 5466
rect 5896 5414 5902 5466
rect 5902 5414 5914 5466
rect 5914 5414 5952 5466
rect 5976 5414 5978 5466
rect 5978 5414 6030 5466
rect 6030 5414 6032 5466
rect 5656 5412 5712 5414
rect 5736 5412 5792 5414
rect 5816 5412 5872 5414
rect 5896 5412 5952 5414
rect 5976 5412 6032 5414
rect 4916 4922 4972 4924
rect 4996 4922 5052 4924
rect 5076 4922 5132 4924
rect 5156 4922 5212 4924
rect 5236 4922 5292 4924
rect 4916 4870 4918 4922
rect 4918 4870 4970 4922
rect 4970 4870 4972 4922
rect 4996 4870 5034 4922
rect 5034 4870 5046 4922
rect 5046 4870 5052 4922
rect 5076 4870 5098 4922
rect 5098 4870 5110 4922
rect 5110 4870 5132 4922
rect 5156 4870 5162 4922
rect 5162 4870 5174 4922
rect 5174 4870 5212 4922
rect 5236 4870 5238 4922
rect 5238 4870 5290 4922
rect 5290 4870 5292 4922
rect 4916 4868 4972 4870
rect 4996 4868 5052 4870
rect 5076 4868 5132 4870
rect 5156 4868 5212 4870
rect 5236 4868 5292 4870
rect 5656 4378 5712 4380
rect 5736 4378 5792 4380
rect 5816 4378 5872 4380
rect 5896 4378 5952 4380
rect 5976 4378 6032 4380
rect 5656 4326 5658 4378
rect 5658 4326 5710 4378
rect 5710 4326 5712 4378
rect 5736 4326 5774 4378
rect 5774 4326 5786 4378
rect 5786 4326 5792 4378
rect 5816 4326 5838 4378
rect 5838 4326 5850 4378
rect 5850 4326 5872 4378
rect 5896 4326 5902 4378
rect 5902 4326 5914 4378
rect 5914 4326 5952 4378
rect 5976 4326 5978 4378
rect 5978 4326 6030 4378
rect 6030 4326 6032 4378
rect 5656 4324 5712 4326
rect 5736 4324 5792 4326
rect 5816 4324 5872 4326
rect 5896 4324 5952 4326
rect 5976 4324 6032 4326
rect 4916 3834 4972 3836
rect 4996 3834 5052 3836
rect 5076 3834 5132 3836
rect 5156 3834 5212 3836
rect 5236 3834 5292 3836
rect 4916 3782 4918 3834
rect 4918 3782 4970 3834
rect 4970 3782 4972 3834
rect 4996 3782 5034 3834
rect 5034 3782 5046 3834
rect 5046 3782 5052 3834
rect 5076 3782 5098 3834
rect 5098 3782 5110 3834
rect 5110 3782 5132 3834
rect 5156 3782 5162 3834
rect 5162 3782 5174 3834
rect 5174 3782 5212 3834
rect 5236 3782 5238 3834
rect 5238 3782 5290 3834
rect 5290 3782 5292 3834
rect 4916 3780 4972 3782
rect 4996 3780 5052 3782
rect 5076 3780 5132 3782
rect 5156 3780 5212 3782
rect 5236 3780 5292 3782
rect 6918 4936 6974 4992
rect 6416 4922 6472 4924
rect 6496 4922 6552 4924
rect 6576 4922 6632 4924
rect 6656 4922 6712 4924
rect 6736 4922 6792 4924
rect 6416 4870 6418 4922
rect 6418 4870 6470 4922
rect 6470 4870 6472 4922
rect 6496 4870 6534 4922
rect 6534 4870 6546 4922
rect 6546 4870 6552 4922
rect 6576 4870 6598 4922
rect 6598 4870 6610 4922
rect 6610 4870 6632 4922
rect 6656 4870 6662 4922
rect 6662 4870 6674 4922
rect 6674 4870 6712 4922
rect 6736 4870 6738 4922
rect 6738 4870 6790 4922
rect 6790 4870 6792 4922
rect 6416 4868 6472 4870
rect 6496 4868 6552 4870
rect 6576 4868 6632 4870
rect 6656 4868 6712 4870
rect 6736 4868 6792 4870
rect 6416 3834 6472 3836
rect 6496 3834 6552 3836
rect 6576 3834 6632 3836
rect 6656 3834 6712 3836
rect 6736 3834 6792 3836
rect 6416 3782 6418 3834
rect 6418 3782 6470 3834
rect 6470 3782 6472 3834
rect 6496 3782 6534 3834
rect 6534 3782 6546 3834
rect 6546 3782 6552 3834
rect 6576 3782 6598 3834
rect 6598 3782 6610 3834
rect 6610 3782 6632 3834
rect 6656 3782 6662 3834
rect 6662 3782 6674 3834
rect 6674 3782 6712 3834
rect 6736 3782 6738 3834
rect 6738 3782 6790 3834
rect 6790 3782 6792 3834
rect 6416 3780 6472 3782
rect 6496 3780 6552 3782
rect 6576 3780 6632 3782
rect 6656 3780 6712 3782
rect 6736 3780 6792 3782
rect 5656 3290 5712 3292
rect 5736 3290 5792 3292
rect 5816 3290 5872 3292
rect 5896 3290 5952 3292
rect 5976 3290 6032 3292
rect 5656 3238 5658 3290
rect 5658 3238 5710 3290
rect 5710 3238 5712 3290
rect 5736 3238 5774 3290
rect 5774 3238 5786 3290
rect 5786 3238 5792 3290
rect 5816 3238 5838 3290
rect 5838 3238 5850 3290
rect 5850 3238 5872 3290
rect 5896 3238 5902 3290
rect 5902 3238 5914 3290
rect 5914 3238 5952 3290
rect 5976 3238 5978 3290
rect 5978 3238 6030 3290
rect 6030 3238 6032 3290
rect 5656 3236 5712 3238
rect 5736 3236 5792 3238
rect 5816 3236 5872 3238
rect 5896 3236 5952 3238
rect 5976 3236 6032 3238
rect 4916 2746 4972 2748
rect 4996 2746 5052 2748
rect 5076 2746 5132 2748
rect 5156 2746 5212 2748
rect 5236 2746 5292 2748
rect 4916 2694 4918 2746
rect 4918 2694 4970 2746
rect 4970 2694 4972 2746
rect 4996 2694 5034 2746
rect 5034 2694 5046 2746
rect 5046 2694 5052 2746
rect 5076 2694 5098 2746
rect 5098 2694 5110 2746
rect 5110 2694 5132 2746
rect 5156 2694 5162 2746
rect 5162 2694 5174 2746
rect 5174 2694 5212 2746
rect 5236 2694 5238 2746
rect 5238 2694 5290 2746
rect 5290 2694 5292 2746
rect 4916 2692 4972 2694
rect 4996 2692 5052 2694
rect 5076 2692 5132 2694
rect 5156 2692 5212 2694
rect 5236 2692 5292 2694
rect 6416 2746 6472 2748
rect 6496 2746 6552 2748
rect 6576 2746 6632 2748
rect 6656 2746 6712 2748
rect 6736 2746 6792 2748
rect 6416 2694 6418 2746
rect 6418 2694 6470 2746
rect 6470 2694 6472 2746
rect 6496 2694 6534 2746
rect 6534 2694 6546 2746
rect 6546 2694 6552 2746
rect 6576 2694 6598 2746
rect 6598 2694 6610 2746
rect 6610 2694 6632 2746
rect 6656 2694 6662 2746
rect 6662 2694 6674 2746
rect 6674 2694 6712 2746
rect 6736 2694 6738 2746
rect 6738 2694 6790 2746
rect 6790 2694 6792 2746
rect 6416 2692 6472 2694
rect 6496 2692 6552 2694
rect 6576 2692 6632 2694
rect 6656 2692 6712 2694
rect 6736 2692 6792 2694
rect 5538 2624 5594 2680
rect 2656 2202 2712 2204
rect 2736 2202 2792 2204
rect 2816 2202 2872 2204
rect 2896 2202 2952 2204
rect 2976 2202 3032 2204
rect 2656 2150 2658 2202
rect 2658 2150 2710 2202
rect 2710 2150 2712 2202
rect 2736 2150 2774 2202
rect 2774 2150 2786 2202
rect 2786 2150 2792 2202
rect 2816 2150 2838 2202
rect 2838 2150 2850 2202
rect 2850 2150 2872 2202
rect 2896 2150 2902 2202
rect 2902 2150 2914 2202
rect 2914 2150 2952 2202
rect 2976 2150 2978 2202
rect 2978 2150 3030 2202
rect 3030 2150 3032 2202
rect 2656 2148 2712 2150
rect 2736 2148 2792 2150
rect 2816 2148 2872 2150
rect 2896 2148 2952 2150
rect 2976 2148 3032 2150
rect 1674 1128 1730 1184
rect 4156 2202 4212 2204
rect 4236 2202 4292 2204
rect 4316 2202 4372 2204
rect 4396 2202 4452 2204
rect 4476 2202 4532 2204
rect 4156 2150 4158 2202
rect 4158 2150 4210 2202
rect 4210 2150 4212 2202
rect 4236 2150 4274 2202
rect 4274 2150 4286 2202
rect 4286 2150 4292 2202
rect 4316 2150 4338 2202
rect 4338 2150 4350 2202
rect 4350 2150 4372 2202
rect 4396 2150 4402 2202
rect 4402 2150 4414 2202
rect 4414 2150 4452 2202
rect 4476 2150 4478 2202
rect 4478 2150 4530 2202
rect 4530 2150 4532 2202
rect 4156 2148 4212 2150
rect 4236 2148 4292 2150
rect 4316 2148 4372 2150
rect 4396 2148 4452 2150
rect 4476 2148 4532 2150
rect 5656 2202 5712 2204
rect 5736 2202 5792 2204
rect 5816 2202 5872 2204
rect 5896 2202 5952 2204
rect 5976 2202 6032 2204
rect 5656 2150 5658 2202
rect 5658 2150 5710 2202
rect 5710 2150 5712 2202
rect 5736 2150 5774 2202
rect 5774 2150 5786 2202
rect 5786 2150 5792 2202
rect 5816 2150 5838 2202
rect 5838 2150 5850 2202
rect 5850 2150 5872 2202
rect 5896 2150 5902 2202
rect 5902 2150 5914 2202
rect 5914 2150 5952 2202
rect 5976 2150 5978 2202
rect 5978 2150 6030 2202
rect 6030 2150 6032 2202
rect 5656 2148 5712 2150
rect 5736 2148 5792 2150
rect 5816 2148 5872 2150
rect 5896 2148 5952 2150
rect 5976 2148 6032 2150
<< metal3 >>
rect 0 8802 800 8832
rect 1393 8802 1459 8805
rect 0 8800 1459 8802
rect 0 8744 1398 8800
rect 1454 8744 1459 8800
rect 0 8742 1459 8744
rect 0 8712 800 8742
rect 1393 8739 1459 8742
rect 2646 7648 3042 7649
rect 2646 7584 2652 7648
rect 2716 7584 2732 7648
rect 2796 7584 2812 7648
rect 2876 7584 2892 7648
rect 2956 7584 2972 7648
rect 3036 7584 3042 7648
rect 2646 7583 3042 7584
rect 4146 7648 4542 7649
rect 4146 7584 4152 7648
rect 4216 7584 4232 7648
rect 4296 7584 4312 7648
rect 4376 7584 4392 7648
rect 4456 7584 4472 7648
rect 4536 7584 4542 7648
rect 4146 7583 4542 7584
rect 5646 7648 6042 7649
rect 5646 7584 5652 7648
rect 5716 7584 5732 7648
rect 5796 7584 5812 7648
rect 5876 7584 5892 7648
rect 5956 7584 5972 7648
rect 6036 7584 6042 7648
rect 5646 7583 6042 7584
rect 1906 7104 2302 7105
rect 1906 7040 1912 7104
rect 1976 7040 1992 7104
rect 2056 7040 2072 7104
rect 2136 7040 2152 7104
rect 2216 7040 2232 7104
rect 2296 7040 2302 7104
rect 1906 7039 2302 7040
rect 3406 7104 3802 7105
rect 3406 7040 3412 7104
rect 3476 7040 3492 7104
rect 3556 7040 3572 7104
rect 3636 7040 3652 7104
rect 3716 7040 3732 7104
rect 3796 7040 3802 7104
rect 3406 7039 3802 7040
rect 4906 7104 5302 7105
rect 4906 7040 4912 7104
rect 4976 7040 4992 7104
rect 5056 7040 5072 7104
rect 5136 7040 5152 7104
rect 5216 7040 5232 7104
rect 5296 7040 5302 7104
rect 4906 7039 5302 7040
rect 6406 7104 6802 7105
rect 6406 7040 6412 7104
rect 6476 7040 6492 7104
rect 6556 7040 6572 7104
rect 6636 7040 6652 7104
rect 6716 7040 6732 7104
rect 6796 7040 6802 7104
rect 6406 7039 6802 7040
rect 0 6898 800 6928
rect 1669 6898 1735 6901
rect 0 6896 1735 6898
rect 0 6840 1674 6896
rect 1730 6840 1735 6896
rect 0 6838 1735 6840
rect 0 6808 800 6838
rect 1669 6835 1735 6838
rect 2646 6560 3042 6561
rect 2646 6496 2652 6560
rect 2716 6496 2732 6560
rect 2796 6496 2812 6560
rect 2876 6496 2892 6560
rect 2956 6496 2972 6560
rect 3036 6496 3042 6560
rect 2646 6495 3042 6496
rect 4146 6560 4542 6561
rect 4146 6496 4152 6560
rect 4216 6496 4232 6560
rect 4296 6496 4312 6560
rect 4376 6496 4392 6560
rect 4456 6496 4472 6560
rect 4536 6496 4542 6560
rect 4146 6495 4542 6496
rect 5646 6560 6042 6561
rect 5646 6496 5652 6560
rect 5716 6496 5732 6560
rect 5796 6496 5812 6560
rect 5876 6496 5892 6560
rect 5956 6496 5972 6560
rect 6036 6496 6042 6560
rect 5646 6495 6042 6496
rect 1906 6016 2302 6017
rect 1906 5952 1912 6016
rect 1976 5952 1992 6016
rect 2056 5952 2072 6016
rect 2136 5952 2152 6016
rect 2216 5952 2232 6016
rect 2296 5952 2302 6016
rect 1906 5951 2302 5952
rect 3406 6016 3802 6017
rect 3406 5952 3412 6016
rect 3476 5952 3492 6016
rect 3556 5952 3572 6016
rect 3636 5952 3652 6016
rect 3716 5952 3732 6016
rect 3796 5952 3802 6016
rect 3406 5951 3802 5952
rect 4906 6016 5302 6017
rect 4906 5952 4912 6016
rect 4976 5952 4992 6016
rect 5056 5952 5072 6016
rect 5136 5952 5152 6016
rect 5216 5952 5232 6016
rect 5296 5952 5302 6016
rect 4906 5951 5302 5952
rect 6406 6016 6802 6017
rect 6406 5952 6412 6016
rect 6476 5952 6492 6016
rect 6556 5952 6572 6016
rect 6636 5952 6652 6016
rect 6716 5952 6732 6016
rect 6796 5952 6802 6016
rect 6406 5951 6802 5952
rect 6085 5676 6151 5677
rect 6085 5674 6132 5676
rect 6040 5672 6132 5674
rect 6040 5616 6090 5672
rect 6040 5614 6132 5616
rect 6085 5612 6132 5614
rect 6196 5612 6202 5676
rect 6085 5611 6151 5612
rect 2646 5472 3042 5473
rect 2646 5408 2652 5472
rect 2716 5408 2732 5472
rect 2796 5408 2812 5472
rect 2876 5408 2892 5472
rect 2956 5408 2972 5472
rect 3036 5408 3042 5472
rect 2646 5407 3042 5408
rect 4146 5472 4542 5473
rect 4146 5408 4152 5472
rect 4216 5408 4232 5472
rect 4296 5408 4312 5472
rect 4376 5408 4392 5472
rect 4456 5408 4472 5472
rect 4536 5408 4542 5472
rect 4146 5407 4542 5408
rect 5646 5472 6042 5473
rect 5646 5408 5652 5472
rect 5716 5408 5732 5472
rect 5796 5408 5812 5472
rect 5876 5408 5892 5472
rect 5956 5408 5972 5472
rect 6036 5408 6042 5472
rect 5646 5407 6042 5408
rect 841 5130 907 5133
rect 798 5128 907 5130
rect 798 5072 846 5128
rect 902 5072 907 5128
rect 798 5067 907 5072
rect 798 5024 858 5067
rect 0 4934 858 5024
rect 6913 4994 6979 4997
rect 7327 4994 8127 5024
rect 6913 4992 8127 4994
rect 6913 4936 6918 4992
rect 6974 4936 8127 4992
rect 6913 4934 8127 4936
rect 0 4904 800 4934
rect 6913 4931 6979 4934
rect 1906 4928 2302 4929
rect 1906 4864 1912 4928
rect 1976 4864 1992 4928
rect 2056 4864 2072 4928
rect 2136 4864 2152 4928
rect 2216 4864 2232 4928
rect 2296 4864 2302 4928
rect 1906 4863 2302 4864
rect 3406 4928 3802 4929
rect 3406 4864 3412 4928
rect 3476 4864 3492 4928
rect 3556 4864 3572 4928
rect 3636 4864 3652 4928
rect 3716 4864 3732 4928
rect 3796 4864 3802 4928
rect 3406 4863 3802 4864
rect 4906 4928 5302 4929
rect 4906 4864 4912 4928
rect 4976 4864 4992 4928
rect 5056 4864 5072 4928
rect 5136 4864 5152 4928
rect 5216 4864 5232 4928
rect 5296 4864 5302 4928
rect 4906 4863 5302 4864
rect 6406 4928 6802 4929
rect 6406 4864 6412 4928
rect 6476 4864 6492 4928
rect 6556 4864 6572 4928
rect 6636 4864 6652 4928
rect 6716 4864 6732 4928
rect 6796 4864 6802 4928
rect 7327 4904 8127 4934
rect 6406 4863 6802 4864
rect 2646 4384 3042 4385
rect 2646 4320 2652 4384
rect 2716 4320 2732 4384
rect 2796 4320 2812 4384
rect 2876 4320 2892 4384
rect 2956 4320 2972 4384
rect 3036 4320 3042 4384
rect 2646 4319 3042 4320
rect 4146 4384 4542 4385
rect 4146 4320 4152 4384
rect 4216 4320 4232 4384
rect 4296 4320 4312 4384
rect 4376 4320 4392 4384
rect 4456 4320 4472 4384
rect 4536 4320 4542 4384
rect 4146 4319 4542 4320
rect 5646 4384 6042 4385
rect 5646 4320 5652 4384
rect 5716 4320 5732 4384
rect 5796 4320 5812 4384
rect 5876 4320 5892 4384
rect 5956 4320 5972 4384
rect 6036 4320 6042 4384
rect 5646 4319 6042 4320
rect 1906 3840 2302 3841
rect 1906 3776 1912 3840
rect 1976 3776 1992 3840
rect 2056 3776 2072 3840
rect 2136 3776 2152 3840
rect 2216 3776 2232 3840
rect 2296 3776 2302 3840
rect 1906 3775 2302 3776
rect 3406 3840 3802 3841
rect 3406 3776 3412 3840
rect 3476 3776 3492 3840
rect 3556 3776 3572 3840
rect 3636 3776 3652 3840
rect 3716 3776 3732 3840
rect 3796 3776 3802 3840
rect 3406 3775 3802 3776
rect 4906 3840 5302 3841
rect 4906 3776 4912 3840
rect 4976 3776 4992 3840
rect 5056 3776 5072 3840
rect 5136 3776 5152 3840
rect 5216 3776 5232 3840
rect 5296 3776 5302 3840
rect 4906 3775 5302 3776
rect 6406 3840 6802 3841
rect 6406 3776 6412 3840
rect 6476 3776 6492 3840
rect 6556 3776 6572 3840
rect 6636 3776 6652 3840
rect 6716 3776 6732 3840
rect 6796 3776 6802 3840
rect 6406 3775 6802 3776
rect 2646 3296 3042 3297
rect 2646 3232 2652 3296
rect 2716 3232 2732 3296
rect 2796 3232 2812 3296
rect 2876 3232 2892 3296
rect 2956 3232 2972 3296
rect 3036 3232 3042 3296
rect 2646 3231 3042 3232
rect 4146 3296 4542 3297
rect 4146 3232 4152 3296
rect 4216 3232 4232 3296
rect 4296 3232 4312 3296
rect 4376 3232 4392 3296
rect 4456 3232 4472 3296
rect 4536 3232 4542 3296
rect 4146 3231 4542 3232
rect 5646 3296 6042 3297
rect 5646 3232 5652 3296
rect 5716 3232 5732 3296
rect 5796 3232 5812 3296
rect 5876 3232 5892 3296
rect 5956 3232 5972 3296
rect 6036 3232 6042 3296
rect 5646 3231 6042 3232
rect 0 3090 800 3120
rect 0 3000 858 3090
rect 798 2957 858 3000
rect 798 2952 907 2957
rect 798 2896 846 2952
rect 902 2896 907 2952
rect 798 2894 907 2896
rect 841 2891 907 2894
rect 1906 2752 2302 2753
rect 1906 2688 1912 2752
rect 1976 2688 1992 2752
rect 2056 2688 2072 2752
rect 2136 2688 2152 2752
rect 2216 2688 2232 2752
rect 2296 2688 2302 2752
rect 1906 2687 2302 2688
rect 3406 2752 3802 2753
rect 3406 2688 3412 2752
rect 3476 2688 3492 2752
rect 3556 2688 3572 2752
rect 3636 2688 3652 2752
rect 3716 2688 3732 2752
rect 3796 2688 3802 2752
rect 3406 2687 3802 2688
rect 4906 2752 5302 2753
rect 4906 2688 4912 2752
rect 4976 2688 4992 2752
rect 5056 2688 5072 2752
rect 5136 2688 5152 2752
rect 5216 2688 5232 2752
rect 5296 2688 5302 2752
rect 4906 2687 5302 2688
rect 6406 2752 6802 2753
rect 6406 2688 6412 2752
rect 6476 2688 6492 2752
rect 6556 2688 6572 2752
rect 6636 2688 6652 2752
rect 6716 2688 6732 2752
rect 6796 2688 6802 2752
rect 6406 2687 6802 2688
rect 5533 2682 5599 2685
rect 6126 2682 6132 2684
rect 5533 2680 6132 2682
rect 5533 2624 5538 2680
rect 5594 2624 6132 2680
rect 5533 2622 6132 2624
rect 5533 2619 5599 2622
rect 6126 2620 6132 2622
rect 6196 2620 6202 2684
rect 2646 2208 3042 2209
rect 2646 2144 2652 2208
rect 2716 2144 2732 2208
rect 2796 2144 2812 2208
rect 2876 2144 2892 2208
rect 2956 2144 2972 2208
rect 3036 2144 3042 2208
rect 2646 2143 3042 2144
rect 4146 2208 4542 2209
rect 4146 2144 4152 2208
rect 4216 2144 4232 2208
rect 4296 2144 4312 2208
rect 4376 2144 4392 2208
rect 4456 2144 4472 2208
rect 4536 2144 4542 2208
rect 4146 2143 4542 2144
rect 5646 2208 6042 2209
rect 5646 2144 5652 2208
rect 5716 2144 5732 2208
rect 5796 2144 5812 2208
rect 5876 2144 5892 2208
rect 5956 2144 5972 2208
rect 6036 2144 6042 2208
rect 5646 2143 6042 2144
rect 0 1186 800 1216
rect 1669 1186 1735 1189
rect 0 1184 1735 1186
rect 0 1128 1674 1184
rect 1730 1128 1735 1184
rect 0 1126 1735 1128
rect 0 1096 800 1126
rect 1669 1123 1735 1126
<< via3 >>
rect 2652 7644 2716 7648
rect 2652 7588 2656 7644
rect 2656 7588 2712 7644
rect 2712 7588 2716 7644
rect 2652 7584 2716 7588
rect 2732 7644 2796 7648
rect 2732 7588 2736 7644
rect 2736 7588 2792 7644
rect 2792 7588 2796 7644
rect 2732 7584 2796 7588
rect 2812 7644 2876 7648
rect 2812 7588 2816 7644
rect 2816 7588 2872 7644
rect 2872 7588 2876 7644
rect 2812 7584 2876 7588
rect 2892 7644 2956 7648
rect 2892 7588 2896 7644
rect 2896 7588 2952 7644
rect 2952 7588 2956 7644
rect 2892 7584 2956 7588
rect 2972 7644 3036 7648
rect 2972 7588 2976 7644
rect 2976 7588 3032 7644
rect 3032 7588 3036 7644
rect 2972 7584 3036 7588
rect 4152 7644 4216 7648
rect 4152 7588 4156 7644
rect 4156 7588 4212 7644
rect 4212 7588 4216 7644
rect 4152 7584 4216 7588
rect 4232 7644 4296 7648
rect 4232 7588 4236 7644
rect 4236 7588 4292 7644
rect 4292 7588 4296 7644
rect 4232 7584 4296 7588
rect 4312 7644 4376 7648
rect 4312 7588 4316 7644
rect 4316 7588 4372 7644
rect 4372 7588 4376 7644
rect 4312 7584 4376 7588
rect 4392 7644 4456 7648
rect 4392 7588 4396 7644
rect 4396 7588 4452 7644
rect 4452 7588 4456 7644
rect 4392 7584 4456 7588
rect 4472 7644 4536 7648
rect 4472 7588 4476 7644
rect 4476 7588 4532 7644
rect 4532 7588 4536 7644
rect 4472 7584 4536 7588
rect 5652 7644 5716 7648
rect 5652 7588 5656 7644
rect 5656 7588 5712 7644
rect 5712 7588 5716 7644
rect 5652 7584 5716 7588
rect 5732 7644 5796 7648
rect 5732 7588 5736 7644
rect 5736 7588 5792 7644
rect 5792 7588 5796 7644
rect 5732 7584 5796 7588
rect 5812 7644 5876 7648
rect 5812 7588 5816 7644
rect 5816 7588 5872 7644
rect 5872 7588 5876 7644
rect 5812 7584 5876 7588
rect 5892 7644 5956 7648
rect 5892 7588 5896 7644
rect 5896 7588 5952 7644
rect 5952 7588 5956 7644
rect 5892 7584 5956 7588
rect 5972 7644 6036 7648
rect 5972 7588 5976 7644
rect 5976 7588 6032 7644
rect 6032 7588 6036 7644
rect 5972 7584 6036 7588
rect 1912 7100 1976 7104
rect 1912 7044 1916 7100
rect 1916 7044 1972 7100
rect 1972 7044 1976 7100
rect 1912 7040 1976 7044
rect 1992 7100 2056 7104
rect 1992 7044 1996 7100
rect 1996 7044 2052 7100
rect 2052 7044 2056 7100
rect 1992 7040 2056 7044
rect 2072 7100 2136 7104
rect 2072 7044 2076 7100
rect 2076 7044 2132 7100
rect 2132 7044 2136 7100
rect 2072 7040 2136 7044
rect 2152 7100 2216 7104
rect 2152 7044 2156 7100
rect 2156 7044 2212 7100
rect 2212 7044 2216 7100
rect 2152 7040 2216 7044
rect 2232 7100 2296 7104
rect 2232 7044 2236 7100
rect 2236 7044 2292 7100
rect 2292 7044 2296 7100
rect 2232 7040 2296 7044
rect 3412 7100 3476 7104
rect 3412 7044 3416 7100
rect 3416 7044 3472 7100
rect 3472 7044 3476 7100
rect 3412 7040 3476 7044
rect 3492 7100 3556 7104
rect 3492 7044 3496 7100
rect 3496 7044 3552 7100
rect 3552 7044 3556 7100
rect 3492 7040 3556 7044
rect 3572 7100 3636 7104
rect 3572 7044 3576 7100
rect 3576 7044 3632 7100
rect 3632 7044 3636 7100
rect 3572 7040 3636 7044
rect 3652 7100 3716 7104
rect 3652 7044 3656 7100
rect 3656 7044 3712 7100
rect 3712 7044 3716 7100
rect 3652 7040 3716 7044
rect 3732 7100 3796 7104
rect 3732 7044 3736 7100
rect 3736 7044 3792 7100
rect 3792 7044 3796 7100
rect 3732 7040 3796 7044
rect 4912 7100 4976 7104
rect 4912 7044 4916 7100
rect 4916 7044 4972 7100
rect 4972 7044 4976 7100
rect 4912 7040 4976 7044
rect 4992 7100 5056 7104
rect 4992 7044 4996 7100
rect 4996 7044 5052 7100
rect 5052 7044 5056 7100
rect 4992 7040 5056 7044
rect 5072 7100 5136 7104
rect 5072 7044 5076 7100
rect 5076 7044 5132 7100
rect 5132 7044 5136 7100
rect 5072 7040 5136 7044
rect 5152 7100 5216 7104
rect 5152 7044 5156 7100
rect 5156 7044 5212 7100
rect 5212 7044 5216 7100
rect 5152 7040 5216 7044
rect 5232 7100 5296 7104
rect 5232 7044 5236 7100
rect 5236 7044 5292 7100
rect 5292 7044 5296 7100
rect 5232 7040 5296 7044
rect 6412 7100 6476 7104
rect 6412 7044 6416 7100
rect 6416 7044 6472 7100
rect 6472 7044 6476 7100
rect 6412 7040 6476 7044
rect 6492 7100 6556 7104
rect 6492 7044 6496 7100
rect 6496 7044 6552 7100
rect 6552 7044 6556 7100
rect 6492 7040 6556 7044
rect 6572 7100 6636 7104
rect 6572 7044 6576 7100
rect 6576 7044 6632 7100
rect 6632 7044 6636 7100
rect 6572 7040 6636 7044
rect 6652 7100 6716 7104
rect 6652 7044 6656 7100
rect 6656 7044 6712 7100
rect 6712 7044 6716 7100
rect 6652 7040 6716 7044
rect 6732 7100 6796 7104
rect 6732 7044 6736 7100
rect 6736 7044 6792 7100
rect 6792 7044 6796 7100
rect 6732 7040 6796 7044
rect 2652 6556 2716 6560
rect 2652 6500 2656 6556
rect 2656 6500 2712 6556
rect 2712 6500 2716 6556
rect 2652 6496 2716 6500
rect 2732 6556 2796 6560
rect 2732 6500 2736 6556
rect 2736 6500 2792 6556
rect 2792 6500 2796 6556
rect 2732 6496 2796 6500
rect 2812 6556 2876 6560
rect 2812 6500 2816 6556
rect 2816 6500 2872 6556
rect 2872 6500 2876 6556
rect 2812 6496 2876 6500
rect 2892 6556 2956 6560
rect 2892 6500 2896 6556
rect 2896 6500 2952 6556
rect 2952 6500 2956 6556
rect 2892 6496 2956 6500
rect 2972 6556 3036 6560
rect 2972 6500 2976 6556
rect 2976 6500 3032 6556
rect 3032 6500 3036 6556
rect 2972 6496 3036 6500
rect 4152 6556 4216 6560
rect 4152 6500 4156 6556
rect 4156 6500 4212 6556
rect 4212 6500 4216 6556
rect 4152 6496 4216 6500
rect 4232 6556 4296 6560
rect 4232 6500 4236 6556
rect 4236 6500 4292 6556
rect 4292 6500 4296 6556
rect 4232 6496 4296 6500
rect 4312 6556 4376 6560
rect 4312 6500 4316 6556
rect 4316 6500 4372 6556
rect 4372 6500 4376 6556
rect 4312 6496 4376 6500
rect 4392 6556 4456 6560
rect 4392 6500 4396 6556
rect 4396 6500 4452 6556
rect 4452 6500 4456 6556
rect 4392 6496 4456 6500
rect 4472 6556 4536 6560
rect 4472 6500 4476 6556
rect 4476 6500 4532 6556
rect 4532 6500 4536 6556
rect 4472 6496 4536 6500
rect 5652 6556 5716 6560
rect 5652 6500 5656 6556
rect 5656 6500 5712 6556
rect 5712 6500 5716 6556
rect 5652 6496 5716 6500
rect 5732 6556 5796 6560
rect 5732 6500 5736 6556
rect 5736 6500 5792 6556
rect 5792 6500 5796 6556
rect 5732 6496 5796 6500
rect 5812 6556 5876 6560
rect 5812 6500 5816 6556
rect 5816 6500 5872 6556
rect 5872 6500 5876 6556
rect 5812 6496 5876 6500
rect 5892 6556 5956 6560
rect 5892 6500 5896 6556
rect 5896 6500 5952 6556
rect 5952 6500 5956 6556
rect 5892 6496 5956 6500
rect 5972 6556 6036 6560
rect 5972 6500 5976 6556
rect 5976 6500 6032 6556
rect 6032 6500 6036 6556
rect 5972 6496 6036 6500
rect 1912 6012 1976 6016
rect 1912 5956 1916 6012
rect 1916 5956 1972 6012
rect 1972 5956 1976 6012
rect 1912 5952 1976 5956
rect 1992 6012 2056 6016
rect 1992 5956 1996 6012
rect 1996 5956 2052 6012
rect 2052 5956 2056 6012
rect 1992 5952 2056 5956
rect 2072 6012 2136 6016
rect 2072 5956 2076 6012
rect 2076 5956 2132 6012
rect 2132 5956 2136 6012
rect 2072 5952 2136 5956
rect 2152 6012 2216 6016
rect 2152 5956 2156 6012
rect 2156 5956 2212 6012
rect 2212 5956 2216 6012
rect 2152 5952 2216 5956
rect 2232 6012 2296 6016
rect 2232 5956 2236 6012
rect 2236 5956 2292 6012
rect 2292 5956 2296 6012
rect 2232 5952 2296 5956
rect 3412 6012 3476 6016
rect 3412 5956 3416 6012
rect 3416 5956 3472 6012
rect 3472 5956 3476 6012
rect 3412 5952 3476 5956
rect 3492 6012 3556 6016
rect 3492 5956 3496 6012
rect 3496 5956 3552 6012
rect 3552 5956 3556 6012
rect 3492 5952 3556 5956
rect 3572 6012 3636 6016
rect 3572 5956 3576 6012
rect 3576 5956 3632 6012
rect 3632 5956 3636 6012
rect 3572 5952 3636 5956
rect 3652 6012 3716 6016
rect 3652 5956 3656 6012
rect 3656 5956 3712 6012
rect 3712 5956 3716 6012
rect 3652 5952 3716 5956
rect 3732 6012 3796 6016
rect 3732 5956 3736 6012
rect 3736 5956 3792 6012
rect 3792 5956 3796 6012
rect 3732 5952 3796 5956
rect 4912 6012 4976 6016
rect 4912 5956 4916 6012
rect 4916 5956 4972 6012
rect 4972 5956 4976 6012
rect 4912 5952 4976 5956
rect 4992 6012 5056 6016
rect 4992 5956 4996 6012
rect 4996 5956 5052 6012
rect 5052 5956 5056 6012
rect 4992 5952 5056 5956
rect 5072 6012 5136 6016
rect 5072 5956 5076 6012
rect 5076 5956 5132 6012
rect 5132 5956 5136 6012
rect 5072 5952 5136 5956
rect 5152 6012 5216 6016
rect 5152 5956 5156 6012
rect 5156 5956 5212 6012
rect 5212 5956 5216 6012
rect 5152 5952 5216 5956
rect 5232 6012 5296 6016
rect 5232 5956 5236 6012
rect 5236 5956 5292 6012
rect 5292 5956 5296 6012
rect 5232 5952 5296 5956
rect 6412 6012 6476 6016
rect 6412 5956 6416 6012
rect 6416 5956 6472 6012
rect 6472 5956 6476 6012
rect 6412 5952 6476 5956
rect 6492 6012 6556 6016
rect 6492 5956 6496 6012
rect 6496 5956 6552 6012
rect 6552 5956 6556 6012
rect 6492 5952 6556 5956
rect 6572 6012 6636 6016
rect 6572 5956 6576 6012
rect 6576 5956 6632 6012
rect 6632 5956 6636 6012
rect 6572 5952 6636 5956
rect 6652 6012 6716 6016
rect 6652 5956 6656 6012
rect 6656 5956 6712 6012
rect 6712 5956 6716 6012
rect 6652 5952 6716 5956
rect 6732 6012 6796 6016
rect 6732 5956 6736 6012
rect 6736 5956 6792 6012
rect 6792 5956 6796 6012
rect 6732 5952 6796 5956
rect 6132 5672 6196 5676
rect 6132 5616 6146 5672
rect 6146 5616 6196 5672
rect 6132 5612 6196 5616
rect 2652 5468 2716 5472
rect 2652 5412 2656 5468
rect 2656 5412 2712 5468
rect 2712 5412 2716 5468
rect 2652 5408 2716 5412
rect 2732 5468 2796 5472
rect 2732 5412 2736 5468
rect 2736 5412 2792 5468
rect 2792 5412 2796 5468
rect 2732 5408 2796 5412
rect 2812 5468 2876 5472
rect 2812 5412 2816 5468
rect 2816 5412 2872 5468
rect 2872 5412 2876 5468
rect 2812 5408 2876 5412
rect 2892 5468 2956 5472
rect 2892 5412 2896 5468
rect 2896 5412 2952 5468
rect 2952 5412 2956 5468
rect 2892 5408 2956 5412
rect 2972 5468 3036 5472
rect 2972 5412 2976 5468
rect 2976 5412 3032 5468
rect 3032 5412 3036 5468
rect 2972 5408 3036 5412
rect 4152 5468 4216 5472
rect 4152 5412 4156 5468
rect 4156 5412 4212 5468
rect 4212 5412 4216 5468
rect 4152 5408 4216 5412
rect 4232 5468 4296 5472
rect 4232 5412 4236 5468
rect 4236 5412 4292 5468
rect 4292 5412 4296 5468
rect 4232 5408 4296 5412
rect 4312 5468 4376 5472
rect 4312 5412 4316 5468
rect 4316 5412 4372 5468
rect 4372 5412 4376 5468
rect 4312 5408 4376 5412
rect 4392 5468 4456 5472
rect 4392 5412 4396 5468
rect 4396 5412 4452 5468
rect 4452 5412 4456 5468
rect 4392 5408 4456 5412
rect 4472 5468 4536 5472
rect 4472 5412 4476 5468
rect 4476 5412 4532 5468
rect 4532 5412 4536 5468
rect 4472 5408 4536 5412
rect 5652 5468 5716 5472
rect 5652 5412 5656 5468
rect 5656 5412 5712 5468
rect 5712 5412 5716 5468
rect 5652 5408 5716 5412
rect 5732 5468 5796 5472
rect 5732 5412 5736 5468
rect 5736 5412 5792 5468
rect 5792 5412 5796 5468
rect 5732 5408 5796 5412
rect 5812 5468 5876 5472
rect 5812 5412 5816 5468
rect 5816 5412 5872 5468
rect 5872 5412 5876 5468
rect 5812 5408 5876 5412
rect 5892 5468 5956 5472
rect 5892 5412 5896 5468
rect 5896 5412 5952 5468
rect 5952 5412 5956 5468
rect 5892 5408 5956 5412
rect 5972 5468 6036 5472
rect 5972 5412 5976 5468
rect 5976 5412 6032 5468
rect 6032 5412 6036 5468
rect 5972 5408 6036 5412
rect 1912 4924 1976 4928
rect 1912 4868 1916 4924
rect 1916 4868 1972 4924
rect 1972 4868 1976 4924
rect 1912 4864 1976 4868
rect 1992 4924 2056 4928
rect 1992 4868 1996 4924
rect 1996 4868 2052 4924
rect 2052 4868 2056 4924
rect 1992 4864 2056 4868
rect 2072 4924 2136 4928
rect 2072 4868 2076 4924
rect 2076 4868 2132 4924
rect 2132 4868 2136 4924
rect 2072 4864 2136 4868
rect 2152 4924 2216 4928
rect 2152 4868 2156 4924
rect 2156 4868 2212 4924
rect 2212 4868 2216 4924
rect 2152 4864 2216 4868
rect 2232 4924 2296 4928
rect 2232 4868 2236 4924
rect 2236 4868 2292 4924
rect 2292 4868 2296 4924
rect 2232 4864 2296 4868
rect 3412 4924 3476 4928
rect 3412 4868 3416 4924
rect 3416 4868 3472 4924
rect 3472 4868 3476 4924
rect 3412 4864 3476 4868
rect 3492 4924 3556 4928
rect 3492 4868 3496 4924
rect 3496 4868 3552 4924
rect 3552 4868 3556 4924
rect 3492 4864 3556 4868
rect 3572 4924 3636 4928
rect 3572 4868 3576 4924
rect 3576 4868 3632 4924
rect 3632 4868 3636 4924
rect 3572 4864 3636 4868
rect 3652 4924 3716 4928
rect 3652 4868 3656 4924
rect 3656 4868 3712 4924
rect 3712 4868 3716 4924
rect 3652 4864 3716 4868
rect 3732 4924 3796 4928
rect 3732 4868 3736 4924
rect 3736 4868 3792 4924
rect 3792 4868 3796 4924
rect 3732 4864 3796 4868
rect 4912 4924 4976 4928
rect 4912 4868 4916 4924
rect 4916 4868 4972 4924
rect 4972 4868 4976 4924
rect 4912 4864 4976 4868
rect 4992 4924 5056 4928
rect 4992 4868 4996 4924
rect 4996 4868 5052 4924
rect 5052 4868 5056 4924
rect 4992 4864 5056 4868
rect 5072 4924 5136 4928
rect 5072 4868 5076 4924
rect 5076 4868 5132 4924
rect 5132 4868 5136 4924
rect 5072 4864 5136 4868
rect 5152 4924 5216 4928
rect 5152 4868 5156 4924
rect 5156 4868 5212 4924
rect 5212 4868 5216 4924
rect 5152 4864 5216 4868
rect 5232 4924 5296 4928
rect 5232 4868 5236 4924
rect 5236 4868 5292 4924
rect 5292 4868 5296 4924
rect 5232 4864 5296 4868
rect 6412 4924 6476 4928
rect 6412 4868 6416 4924
rect 6416 4868 6472 4924
rect 6472 4868 6476 4924
rect 6412 4864 6476 4868
rect 6492 4924 6556 4928
rect 6492 4868 6496 4924
rect 6496 4868 6552 4924
rect 6552 4868 6556 4924
rect 6492 4864 6556 4868
rect 6572 4924 6636 4928
rect 6572 4868 6576 4924
rect 6576 4868 6632 4924
rect 6632 4868 6636 4924
rect 6572 4864 6636 4868
rect 6652 4924 6716 4928
rect 6652 4868 6656 4924
rect 6656 4868 6712 4924
rect 6712 4868 6716 4924
rect 6652 4864 6716 4868
rect 6732 4924 6796 4928
rect 6732 4868 6736 4924
rect 6736 4868 6792 4924
rect 6792 4868 6796 4924
rect 6732 4864 6796 4868
rect 2652 4380 2716 4384
rect 2652 4324 2656 4380
rect 2656 4324 2712 4380
rect 2712 4324 2716 4380
rect 2652 4320 2716 4324
rect 2732 4380 2796 4384
rect 2732 4324 2736 4380
rect 2736 4324 2792 4380
rect 2792 4324 2796 4380
rect 2732 4320 2796 4324
rect 2812 4380 2876 4384
rect 2812 4324 2816 4380
rect 2816 4324 2872 4380
rect 2872 4324 2876 4380
rect 2812 4320 2876 4324
rect 2892 4380 2956 4384
rect 2892 4324 2896 4380
rect 2896 4324 2952 4380
rect 2952 4324 2956 4380
rect 2892 4320 2956 4324
rect 2972 4380 3036 4384
rect 2972 4324 2976 4380
rect 2976 4324 3032 4380
rect 3032 4324 3036 4380
rect 2972 4320 3036 4324
rect 4152 4380 4216 4384
rect 4152 4324 4156 4380
rect 4156 4324 4212 4380
rect 4212 4324 4216 4380
rect 4152 4320 4216 4324
rect 4232 4380 4296 4384
rect 4232 4324 4236 4380
rect 4236 4324 4292 4380
rect 4292 4324 4296 4380
rect 4232 4320 4296 4324
rect 4312 4380 4376 4384
rect 4312 4324 4316 4380
rect 4316 4324 4372 4380
rect 4372 4324 4376 4380
rect 4312 4320 4376 4324
rect 4392 4380 4456 4384
rect 4392 4324 4396 4380
rect 4396 4324 4452 4380
rect 4452 4324 4456 4380
rect 4392 4320 4456 4324
rect 4472 4380 4536 4384
rect 4472 4324 4476 4380
rect 4476 4324 4532 4380
rect 4532 4324 4536 4380
rect 4472 4320 4536 4324
rect 5652 4380 5716 4384
rect 5652 4324 5656 4380
rect 5656 4324 5712 4380
rect 5712 4324 5716 4380
rect 5652 4320 5716 4324
rect 5732 4380 5796 4384
rect 5732 4324 5736 4380
rect 5736 4324 5792 4380
rect 5792 4324 5796 4380
rect 5732 4320 5796 4324
rect 5812 4380 5876 4384
rect 5812 4324 5816 4380
rect 5816 4324 5872 4380
rect 5872 4324 5876 4380
rect 5812 4320 5876 4324
rect 5892 4380 5956 4384
rect 5892 4324 5896 4380
rect 5896 4324 5952 4380
rect 5952 4324 5956 4380
rect 5892 4320 5956 4324
rect 5972 4380 6036 4384
rect 5972 4324 5976 4380
rect 5976 4324 6032 4380
rect 6032 4324 6036 4380
rect 5972 4320 6036 4324
rect 1912 3836 1976 3840
rect 1912 3780 1916 3836
rect 1916 3780 1972 3836
rect 1972 3780 1976 3836
rect 1912 3776 1976 3780
rect 1992 3836 2056 3840
rect 1992 3780 1996 3836
rect 1996 3780 2052 3836
rect 2052 3780 2056 3836
rect 1992 3776 2056 3780
rect 2072 3836 2136 3840
rect 2072 3780 2076 3836
rect 2076 3780 2132 3836
rect 2132 3780 2136 3836
rect 2072 3776 2136 3780
rect 2152 3836 2216 3840
rect 2152 3780 2156 3836
rect 2156 3780 2212 3836
rect 2212 3780 2216 3836
rect 2152 3776 2216 3780
rect 2232 3836 2296 3840
rect 2232 3780 2236 3836
rect 2236 3780 2292 3836
rect 2292 3780 2296 3836
rect 2232 3776 2296 3780
rect 3412 3836 3476 3840
rect 3412 3780 3416 3836
rect 3416 3780 3472 3836
rect 3472 3780 3476 3836
rect 3412 3776 3476 3780
rect 3492 3836 3556 3840
rect 3492 3780 3496 3836
rect 3496 3780 3552 3836
rect 3552 3780 3556 3836
rect 3492 3776 3556 3780
rect 3572 3836 3636 3840
rect 3572 3780 3576 3836
rect 3576 3780 3632 3836
rect 3632 3780 3636 3836
rect 3572 3776 3636 3780
rect 3652 3836 3716 3840
rect 3652 3780 3656 3836
rect 3656 3780 3712 3836
rect 3712 3780 3716 3836
rect 3652 3776 3716 3780
rect 3732 3836 3796 3840
rect 3732 3780 3736 3836
rect 3736 3780 3792 3836
rect 3792 3780 3796 3836
rect 3732 3776 3796 3780
rect 4912 3836 4976 3840
rect 4912 3780 4916 3836
rect 4916 3780 4972 3836
rect 4972 3780 4976 3836
rect 4912 3776 4976 3780
rect 4992 3836 5056 3840
rect 4992 3780 4996 3836
rect 4996 3780 5052 3836
rect 5052 3780 5056 3836
rect 4992 3776 5056 3780
rect 5072 3836 5136 3840
rect 5072 3780 5076 3836
rect 5076 3780 5132 3836
rect 5132 3780 5136 3836
rect 5072 3776 5136 3780
rect 5152 3836 5216 3840
rect 5152 3780 5156 3836
rect 5156 3780 5212 3836
rect 5212 3780 5216 3836
rect 5152 3776 5216 3780
rect 5232 3836 5296 3840
rect 5232 3780 5236 3836
rect 5236 3780 5292 3836
rect 5292 3780 5296 3836
rect 5232 3776 5296 3780
rect 6412 3836 6476 3840
rect 6412 3780 6416 3836
rect 6416 3780 6472 3836
rect 6472 3780 6476 3836
rect 6412 3776 6476 3780
rect 6492 3836 6556 3840
rect 6492 3780 6496 3836
rect 6496 3780 6552 3836
rect 6552 3780 6556 3836
rect 6492 3776 6556 3780
rect 6572 3836 6636 3840
rect 6572 3780 6576 3836
rect 6576 3780 6632 3836
rect 6632 3780 6636 3836
rect 6572 3776 6636 3780
rect 6652 3836 6716 3840
rect 6652 3780 6656 3836
rect 6656 3780 6712 3836
rect 6712 3780 6716 3836
rect 6652 3776 6716 3780
rect 6732 3836 6796 3840
rect 6732 3780 6736 3836
rect 6736 3780 6792 3836
rect 6792 3780 6796 3836
rect 6732 3776 6796 3780
rect 2652 3292 2716 3296
rect 2652 3236 2656 3292
rect 2656 3236 2712 3292
rect 2712 3236 2716 3292
rect 2652 3232 2716 3236
rect 2732 3292 2796 3296
rect 2732 3236 2736 3292
rect 2736 3236 2792 3292
rect 2792 3236 2796 3292
rect 2732 3232 2796 3236
rect 2812 3292 2876 3296
rect 2812 3236 2816 3292
rect 2816 3236 2872 3292
rect 2872 3236 2876 3292
rect 2812 3232 2876 3236
rect 2892 3292 2956 3296
rect 2892 3236 2896 3292
rect 2896 3236 2952 3292
rect 2952 3236 2956 3292
rect 2892 3232 2956 3236
rect 2972 3292 3036 3296
rect 2972 3236 2976 3292
rect 2976 3236 3032 3292
rect 3032 3236 3036 3292
rect 2972 3232 3036 3236
rect 4152 3292 4216 3296
rect 4152 3236 4156 3292
rect 4156 3236 4212 3292
rect 4212 3236 4216 3292
rect 4152 3232 4216 3236
rect 4232 3292 4296 3296
rect 4232 3236 4236 3292
rect 4236 3236 4292 3292
rect 4292 3236 4296 3292
rect 4232 3232 4296 3236
rect 4312 3292 4376 3296
rect 4312 3236 4316 3292
rect 4316 3236 4372 3292
rect 4372 3236 4376 3292
rect 4312 3232 4376 3236
rect 4392 3292 4456 3296
rect 4392 3236 4396 3292
rect 4396 3236 4452 3292
rect 4452 3236 4456 3292
rect 4392 3232 4456 3236
rect 4472 3292 4536 3296
rect 4472 3236 4476 3292
rect 4476 3236 4532 3292
rect 4532 3236 4536 3292
rect 4472 3232 4536 3236
rect 5652 3292 5716 3296
rect 5652 3236 5656 3292
rect 5656 3236 5712 3292
rect 5712 3236 5716 3292
rect 5652 3232 5716 3236
rect 5732 3292 5796 3296
rect 5732 3236 5736 3292
rect 5736 3236 5792 3292
rect 5792 3236 5796 3292
rect 5732 3232 5796 3236
rect 5812 3292 5876 3296
rect 5812 3236 5816 3292
rect 5816 3236 5872 3292
rect 5872 3236 5876 3292
rect 5812 3232 5876 3236
rect 5892 3292 5956 3296
rect 5892 3236 5896 3292
rect 5896 3236 5952 3292
rect 5952 3236 5956 3292
rect 5892 3232 5956 3236
rect 5972 3292 6036 3296
rect 5972 3236 5976 3292
rect 5976 3236 6032 3292
rect 6032 3236 6036 3292
rect 5972 3232 6036 3236
rect 1912 2748 1976 2752
rect 1912 2692 1916 2748
rect 1916 2692 1972 2748
rect 1972 2692 1976 2748
rect 1912 2688 1976 2692
rect 1992 2748 2056 2752
rect 1992 2692 1996 2748
rect 1996 2692 2052 2748
rect 2052 2692 2056 2748
rect 1992 2688 2056 2692
rect 2072 2748 2136 2752
rect 2072 2692 2076 2748
rect 2076 2692 2132 2748
rect 2132 2692 2136 2748
rect 2072 2688 2136 2692
rect 2152 2748 2216 2752
rect 2152 2692 2156 2748
rect 2156 2692 2212 2748
rect 2212 2692 2216 2748
rect 2152 2688 2216 2692
rect 2232 2748 2296 2752
rect 2232 2692 2236 2748
rect 2236 2692 2292 2748
rect 2292 2692 2296 2748
rect 2232 2688 2296 2692
rect 3412 2748 3476 2752
rect 3412 2692 3416 2748
rect 3416 2692 3472 2748
rect 3472 2692 3476 2748
rect 3412 2688 3476 2692
rect 3492 2748 3556 2752
rect 3492 2692 3496 2748
rect 3496 2692 3552 2748
rect 3552 2692 3556 2748
rect 3492 2688 3556 2692
rect 3572 2748 3636 2752
rect 3572 2692 3576 2748
rect 3576 2692 3632 2748
rect 3632 2692 3636 2748
rect 3572 2688 3636 2692
rect 3652 2748 3716 2752
rect 3652 2692 3656 2748
rect 3656 2692 3712 2748
rect 3712 2692 3716 2748
rect 3652 2688 3716 2692
rect 3732 2748 3796 2752
rect 3732 2692 3736 2748
rect 3736 2692 3792 2748
rect 3792 2692 3796 2748
rect 3732 2688 3796 2692
rect 4912 2748 4976 2752
rect 4912 2692 4916 2748
rect 4916 2692 4972 2748
rect 4972 2692 4976 2748
rect 4912 2688 4976 2692
rect 4992 2748 5056 2752
rect 4992 2692 4996 2748
rect 4996 2692 5052 2748
rect 5052 2692 5056 2748
rect 4992 2688 5056 2692
rect 5072 2748 5136 2752
rect 5072 2692 5076 2748
rect 5076 2692 5132 2748
rect 5132 2692 5136 2748
rect 5072 2688 5136 2692
rect 5152 2748 5216 2752
rect 5152 2692 5156 2748
rect 5156 2692 5212 2748
rect 5212 2692 5216 2748
rect 5152 2688 5216 2692
rect 5232 2748 5296 2752
rect 5232 2692 5236 2748
rect 5236 2692 5292 2748
rect 5292 2692 5296 2748
rect 5232 2688 5296 2692
rect 6412 2748 6476 2752
rect 6412 2692 6416 2748
rect 6416 2692 6472 2748
rect 6472 2692 6476 2748
rect 6412 2688 6476 2692
rect 6492 2748 6556 2752
rect 6492 2692 6496 2748
rect 6496 2692 6552 2748
rect 6552 2692 6556 2748
rect 6492 2688 6556 2692
rect 6572 2748 6636 2752
rect 6572 2692 6576 2748
rect 6576 2692 6632 2748
rect 6632 2692 6636 2748
rect 6572 2688 6636 2692
rect 6652 2748 6716 2752
rect 6652 2692 6656 2748
rect 6656 2692 6712 2748
rect 6712 2692 6716 2748
rect 6652 2688 6716 2692
rect 6732 2748 6796 2752
rect 6732 2692 6736 2748
rect 6736 2692 6792 2748
rect 6792 2692 6796 2748
rect 6732 2688 6796 2692
rect 6132 2620 6196 2684
rect 2652 2204 2716 2208
rect 2652 2148 2656 2204
rect 2656 2148 2712 2204
rect 2712 2148 2716 2204
rect 2652 2144 2716 2148
rect 2732 2204 2796 2208
rect 2732 2148 2736 2204
rect 2736 2148 2792 2204
rect 2792 2148 2796 2204
rect 2732 2144 2796 2148
rect 2812 2204 2876 2208
rect 2812 2148 2816 2204
rect 2816 2148 2872 2204
rect 2872 2148 2876 2204
rect 2812 2144 2876 2148
rect 2892 2204 2956 2208
rect 2892 2148 2896 2204
rect 2896 2148 2952 2204
rect 2952 2148 2956 2204
rect 2892 2144 2956 2148
rect 2972 2204 3036 2208
rect 2972 2148 2976 2204
rect 2976 2148 3032 2204
rect 3032 2148 3036 2204
rect 2972 2144 3036 2148
rect 4152 2204 4216 2208
rect 4152 2148 4156 2204
rect 4156 2148 4212 2204
rect 4212 2148 4216 2204
rect 4152 2144 4216 2148
rect 4232 2204 4296 2208
rect 4232 2148 4236 2204
rect 4236 2148 4292 2204
rect 4292 2148 4296 2204
rect 4232 2144 4296 2148
rect 4312 2204 4376 2208
rect 4312 2148 4316 2204
rect 4316 2148 4372 2204
rect 4372 2148 4376 2204
rect 4312 2144 4376 2148
rect 4392 2204 4456 2208
rect 4392 2148 4396 2204
rect 4396 2148 4452 2204
rect 4452 2148 4456 2204
rect 4392 2144 4456 2148
rect 4472 2204 4536 2208
rect 4472 2148 4476 2204
rect 4476 2148 4532 2204
rect 4532 2148 4536 2204
rect 4472 2144 4536 2148
rect 5652 2204 5716 2208
rect 5652 2148 5656 2204
rect 5656 2148 5712 2204
rect 5712 2148 5716 2204
rect 5652 2144 5716 2148
rect 5732 2204 5796 2208
rect 5732 2148 5736 2204
rect 5736 2148 5792 2204
rect 5792 2148 5796 2204
rect 5732 2144 5796 2148
rect 5812 2204 5876 2208
rect 5812 2148 5816 2204
rect 5816 2148 5872 2204
rect 5872 2148 5876 2204
rect 5812 2144 5876 2148
rect 5892 2204 5956 2208
rect 5892 2148 5896 2204
rect 5896 2148 5952 2204
rect 5952 2148 5956 2204
rect 5892 2144 5956 2148
rect 5972 2204 6036 2208
rect 5972 2148 5976 2204
rect 5976 2148 6032 2204
rect 6032 2148 6036 2204
rect 5972 2144 6036 2148
<< metal4 >>
rect 1904 7104 2304 7664
rect 1904 7040 1912 7104
rect 1976 7040 1992 7104
rect 2056 7040 2072 7104
rect 2136 7040 2152 7104
rect 2216 7040 2232 7104
rect 2296 7040 2304 7104
rect 1904 6016 2304 7040
rect 1904 5952 1912 6016
rect 1976 5952 1992 6016
rect 2056 5952 2072 6016
rect 2136 5952 2152 6016
rect 2216 5952 2232 6016
rect 2296 5952 2304 6016
rect 1904 4928 2304 5952
rect 1904 4864 1912 4928
rect 1976 4864 1992 4928
rect 2056 4864 2072 4928
rect 2136 4864 2152 4928
rect 2216 4864 2232 4928
rect 2296 4864 2304 4928
rect 1904 3840 2304 4864
rect 1904 3776 1912 3840
rect 1976 3776 1992 3840
rect 2056 3776 2072 3840
rect 2136 3776 2152 3840
rect 2216 3776 2232 3840
rect 2296 3776 2304 3840
rect 1904 2752 2304 3776
rect 1904 2688 1912 2752
rect 1976 2688 1992 2752
rect 2056 2688 2072 2752
rect 2136 2688 2152 2752
rect 2216 2688 2232 2752
rect 2296 2688 2304 2752
rect 1904 2128 2304 2688
rect 2644 7648 3044 7664
rect 2644 7584 2652 7648
rect 2716 7584 2732 7648
rect 2796 7584 2812 7648
rect 2876 7584 2892 7648
rect 2956 7584 2972 7648
rect 3036 7584 3044 7648
rect 2644 6560 3044 7584
rect 2644 6496 2652 6560
rect 2716 6496 2732 6560
rect 2796 6496 2812 6560
rect 2876 6496 2892 6560
rect 2956 6496 2972 6560
rect 3036 6496 3044 6560
rect 2644 5472 3044 6496
rect 2644 5408 2652 5472
rect 2716 5408 2732 5472
rect 2796 5408 2812 5472
rect 2876 5408 2892 5472
rect 2956 5408 2972 5472
rect 3036 5408 3044 5472
rect 2644 4384 3044 5408
rect 2644 4320 2652 4384
rect 2716 4320 2732 4384
rect 2796 4320 2812 4384
rect 2876 4320 2892 4384
rect 2956 4320 2972 4384
rect 3036 4320 3044 4384
rect 2644 3296 3044 4320
rect 2644 3232 2652 3296
rect 2716 3232 2732 3296
rect 2796 3232 2812 3296
rect 2876 3232 2892 3296
rect 2956 3232 2972 3296
rect 3036 3232 3044 3296
rect 2644 2208 3044 3232
rect 2644 2144 2652 2208
rect 2716 2144 2732 2208
rect 2796 2144 2812 2208
rect 2876 2144 2892 2208
rect 2956 2144 2972 2208
rect 3036 2144 3044 2208
rect 2644 2128 3044 2144
rect 3404 7104 3804 7664
rect 3404 7040 3412 7104
rect 3476 7040 3492 7104
rect 3556 7040 3572 7104
rect 3636 7040 3652 7104
rect 3716 7040 3732 7104
rect 3796 7040 3804 7104
rect 3404 6016 3804 7040
rect 3404 5952 3412 6016
rect 3476 5952 3492 6016
rect 3556 5952 3572 6016
rect 3636 5952 3652 6016
rect 3716 5952 3732 6016
rect 3796 5952 3804 6016
rect 3404 4928 3804 5952
rect 3404 4864 3412 4928
rect 3476 4864 3492 4928
rect 3556 4864 3572 4928
rect 3636 4864 3652 4928
rect 3716 4864 3732 4928
rect 3796 4864 3804 4928
rect 3404 3840 3804 4864
rect 3404 3776 3412 3840
rect 3476 3776 3492 3840
rect 3556 3776 3572 3840
rect 3636 3776 3652 3840
rect 3716 3776 3732 3840
rect 3796 3776 3804 3840
rect 3404 2752 3804 3776
rect 3404 2688 3412 2752
rect 3476 2688 3492 2752
rect 3556 2688 3572 2752
rect 3636 2688 3652 2752
rect 3716 2688 3732 2752
rect 3796 2688 3804 2752
rect 3404 2128 3804 2688
rect 4144 7648 4544 7664
rect 4144 7584 4152 7648
rect 4216 7584 4232 7648
rect 4296 7584 4312 7648
rect 4376 7584 4392 7648
rect 4456 7584 4472 7648
rect 4536 7584 4544 7648
rect 4144 6560 4544 7584
rect 4144 6496 4152 6560
rect 4216 6496 4232 6560
rect 4296 6496 4312 6560
rect 4376 6496 4392 6560
rect 4456 6496 4472 6560
rect 4536 6496 4544 6560
rect 4144 5472 4544 6496
rect 4144 5408 4152 5472
rect 4216 5408 4232 5472
rect 4296 5408 4312 5472
rect 4376 5408 4392 5472
rect 4456 5408 4472 5472
rect 4536 5408 4544 5472
rect 4144 4384 4544 5408
rect 4144 4320 4152 4384
rect 4216 4320 4232 4384
rect 4296 4320 4312 4384
rect 4376 4320 4392 4384
rect 4456 4320 4472 4384
rect 4536 4320 4544 4384
rect 4144 3296 4544 4320
rect 4144 3232 4152 3296
rect 4216 3232 4232 3296
rect 4296 3232 4312 3296
rect 4376 3232 4392 3296
rect 4456 3232 4472 3296
rect 4536 3232 4544 3296
rect 4144 2208 4544 3232
rect 4144 2144 4152 2208
rect 4216 2144 4232 2208
rect 4296 2144 4312 2208
rect 4376 2144 4392 2208
rect 4456 2144 4472 2208
rect 4536 2144 4544 2208
rect 4144 2128 4544 2144
rect 4904 7104 5304 7664
rect 4904 7040 4912 7104
rect 4976 7040 4992 7104
rect 5056 7040 5072 7104
rect 5136 7040 5152 7104
rect 5216 7040 5232 7104
rect 5296 7040 5304 7104
rect 4904 6016 5304 7040
rect 4904 5952 4912 6016
rect 4976 5952 4992 6016
rect 5056 5952 5072 6016
rect 5136 5952 5152 6016
rect 5216 5952 5232 6016
rect 5296 5952 5304 6016
rect 4904 4928 5304 5952
rect 4904 4864 4912 4928
rect 4976 4864 4992 4928
rect 5056 4864 5072 4928
rect 5136 4864 5152 4928
rect 5216 4864 5232 4928
rect 5296 4864 5304 4928
rect 4904 3840 5304 4864
rect 4904 3776 4912 3840
rect 4976 3776 4992 3840
rect 5056 3776 5072 3840
rect 5136 3776 5152 3840
rect 5216 3776 5232 3840
rect 5296 3776 5304 3840
rect 4904 2752 5304 3776
rect 4904 2688 4912 2752
rect 4976 2688 4992 2752
rect 5056 2688 5072 2752
rect 5136 2688 5152 2752
rect 5216 2688 5232 2752
rect 5296 2688 5304 2752
rect 4904 2128 5304 2688
rect 5644 7648 6044 7664
rect 5644 7584 5652 7648
rect 5716 7584 5732 7648
rect 5796 7584 5812 7648
rect 5876 7584 5892 7648
rect 5956 7584 5972 7648
rect 6036 7584 6044 7648
rect 5644 6560 6044 7584
rect 5644 6496 5652 6560
rect 5716 6496 5732 6560
rect 5796 6496 5812 6560
rect 5876 6496 5892 6560
rect 5956 6496 5972 6560
rect 6036 6496 6044 6560
rect 5644 5472 6044 6496
rect 6404 7104 6804 7664
rect 6404 7040 6412 7104
rect 6476 7040 6492 7104
rect 6556 7040 6572 7104
rect 6636 7040 6652 7104
rect 6716 7040 6732 7104
rect 6796 7040 6804 7104
rect 6404 6016 6804 7040
rect 6404 5952 6412 6016
rect 6476 5952 6492 6016
rect 6556 5952 6572 6016
rect 6636 5952 6652 6016
rect 6716 5952 6732 6016
rect 6796 5952 6804 6016
rect 6131 5676 6197 5677
rect 6131 5612 6132 5676
rect 6196 5612 6197 5676
rect 6131 5611 6197 5612
rect 5644 5408 5652 5472
rect 5716 5408 5732 5472
rect 5796 5408 5812 5472
rect 5876 5408 5892 5472
rect 5956 5408 5972 5472
rect 6036 5408 6044 5472
rect 5644 4384 6044 5408
rect 5644 4320 5652 4384
rect 5716 4320 5732 4384
rect 5796 4320 5812 4384
rect 5876 4320 5892 4384
rect 5956 4320 5972 4384
rect 6036 4320 6044 4384
rect 5644 3296 6044 4320
rect 5644 3232 5652 3296
rect 5716 3232 5732 3296
rect 5796 3232 5812 3296
rect 5876 3232 5892 3296
rect 5956 3232 5972 3296
rect 6036 3232 6044 3296
rect 5644 2208 6044 3232
rect 6134 2685 6194 5611
rect 6404 4928 6804 5952
rect 6404 4864 6412 4928
rect 6476 4864 6492 4928
rect 6556 4864 6572 4928
rect 6636 4864 6652 4928
rect 6716 4864 6732 4928
rect 6796 4864 6804 4928
rect 6404 3840 6804 4864
rect 6404 3776 6412 3840
rect 6476 3776 6492 3840
rect 6556 3776 6572 3840
rect 6636 3776 6652 3840
rect 6716 3776 6732 3840
rect 6796 3776 6804 3840
rect 6404 2752 6804 3776
rect 6404 2688 6412 2752
rect 6476 2688 6492 2752
rect 6556 2688 6572 2752
rect 6636 2688 6652 2752
rect 6716 2688 6732 2752
rect 6796 2688 6804 2752
rect 6131 2684 6197 2685
rect 6131 2620 6132 2684
rect 6196 2620 6197 2684
rect 6131 2619 6197 2620
rect 5644 2144 5652 2208
rect 5716 2144 5732 2208
rect 5796 2144 5812 2208
rect 5876 2144 5892 2208
rect 5956 2144 5972 2208
rect 6036 2144 6044 2208
rect 5644 2128 6044 2144
rect 6404 2128 6804 2688
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CLK ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 5612 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CLK
timestamp 1704896540
transform -1 0 3220 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CLK
timestamp 1704896540
transform 1 0 4876 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_23 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3220 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_49 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_57 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_9
timestamp 1704896540
transform 1 0 1932 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_37 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4508 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_49
timestamp 1704896540
transform 1 0 5612 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1704896540
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_57
timestamp 1704896540
transform 1 0 6348 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_3
timestamp 1704896540
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_52 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5888 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_60
timestamp 1704896540
transform 1 0 6624 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_3
timestamp 1704896540
transform 1 0 1380 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_11
timestamp 1704896540
transform 1 0 2116 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1704896540
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1704896540
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1704896540
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_57
timestamp 1704896540
transform 1 0 6348 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_3
timestamp 1704896540
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_55
timestamp 1704896540
transform 1 0 6164 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_6
timestamp 1704896540
transform 1 0 1656 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_18
timestamp 1704896540
transform 1 0 2760 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_48
timestamp 1704896540
transform 1 0 5520 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_57
timestamp 1704896540
transform 1 0 6348 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_3
timestamp 1704896540
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_52
timestamp 1704896540
transform 1 0 5888 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_60
timestamp 1704896540
transform 1 0 6624 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1704896540
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_41
timestamp 1704896540
transform 1 0 4876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_53 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_57
timestamp 1704896540
transform 1 0 6348 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1704896540
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1704896540
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1704896540
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1704896540
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_9
timestamp 1704896540
transform 1 0 1932 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_14
timestamp 1704896540
transform 1 0 2392 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_26
timestamp 1704896540
transform 1 0 3496 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_29
timestamp 1704896540
transform 1 0 3772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_41
timestamp 1704896540
transform 1 0 4876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_53
timestamp 1704896540
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_57
timestamp 1704896540
transform 1 0 6348 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input1 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 3680 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input2 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2024 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1704896540
transform -1 0 6716 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output4
timestamp 1704896540
transform -1 0 1932 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output5
timestamp 1704896540
transform -1 0 1656 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output6
timestamp 1704896540
transform -1 0 1656 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output7
timestamp 1704896540
transform -1 0 1932 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output8
timestamp 1704896540
transform -1 0 1656 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_10
timestamp 1704896540
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1704896540
transform -1 0 6992 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_11
timestamp 1704896540
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1704896540
transform -1 0 6992 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_12
timestamp 1704896540
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1704896540
transform -1 0 6992 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_13
timestamp 1704896540
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1704896540
transform -1 0 6992 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_14
timestamp 1704896540
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1704896540
transform -1 0 6992 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_15
timestamp 1704896540
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1704896540
transform -1 0 6992 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_16
timestamp 1704896540
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1704896540
transform -1 0 6992 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_17
timestamp 1704896540
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1704896540
transform -1 0 6992 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_18
timestamp 1704896540
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1704896540
transform -1 0 6992 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_19
timestamp 1704896540
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1704896540
transform -1 0 6992 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_20 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_21
timestamp 1704896540
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_22
timestamp 1704896540
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_23
timestamp 1704896540
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_24
timestamp 1704896540
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_25
timestamp 1704896540
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_26
timestamp 1704896540
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_27
timestamp 1704896540
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_28
timestamp 1704896540
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_29
timestamp 1704896540
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_30
timestamp 1704896540
transform 1 0 3680 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_31
timestamp 1704896540
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__dfrbp_1  x1 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1564 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrbp_1  x2
timestamp 1704896540
transform 1 0 1564 0 1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfsbp_1  x3 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 5888 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrbp_1  x4
timestamp 1704896540
transform 1 0 1564 0 1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrbp_1  x5
timestamp 1704896540
transform -1 0 5888 0 1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfbbp_1  x6 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 4508 0 -1 3264
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbp_1  x7
timestamp 1704896540
transform -1 0 6164 0 1 4352
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbp_1  x8
timestamp 1704896540
transform -1 0 4692 0 -1 4352
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbp_1  x9
timestamp 1704896540
transform -1 0 5520 0 -1 5440
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbp_1  x10
timestamp 1704896540
transform 1 0 2484 0 -1 6528
box -38 -48 2430 592
<< labels >>
flabel metal2 s 5998 9471 6054 10271 0 FreeSans 224 90 0 0 CLK
port 0 nsew signal input
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 D0
port 1 nsew signal output
flabel metal3 s 0 4904 800 5024 0 FreeSans 480 0 0 0 D1
port 2 nsew signal output
flabel metal3 s 0 3000 800 3120 0 FreeSans 480 0 0 0 D2
port 3 nsew signal output
flabel metal3 s 0 1096 800 1216 0 FreeSans 480 0 0 0 D3
port 4 nsew signal output
flabel metal3 s 0 8712 800 8832 0 FreeSans 480 0 0 0 EOC
port 5 nsew signal output
flabel metal2 s 3974 0 4030 800 0 FreeSans 224 90 0 0 GND
port 6 nsew signal input
flabel metal2 s 1950 9471 2006 10271 0 FreeSans 224 90 0 0 NRST
port 7 nsew signal input
flabel metal4 s 2644 2128 3044 7664 0 FreeSans 1920 90 0 0 VGND
port 8 nsew ground bidirectional
flabel metal4 s 4144 2128 4544 7664 0 FreeSans 1920 90 0 0 VGND
port 8 nsew ground bidirectional
flabel metal4 s 5644 2128 6044 7664 0 FreeSans 1920 90 0 0 VGND
port 8 nsew ground bidirectional
flabel metal4 s 1904 2128 2304 7664 0 FreeSans 1920 90 0 0 VPWR
port 9 nsew power bidirectional
flabel metal4 s 3404 2128 3804 7664 0 FreeSans 1920 90 0 0 VPWR
port 9 nsew power bidirectional
flabel metal4 s 4904 2128 5304 7664 0 FreeSans 1920 90 0 0 VPWR
port 9 nsew power bidirectional
flabel metal4 s 6404 2128 6804 7664 0 FreeSans 1920 90 0 0 VPWR
port 9 nsew power bidirectional
flabel metal3 s 7327 4904 8127 5024 0 FreeSans 480 0 0 0 Vcomp
port 10 nsew signal input
rlabel metal1 4048 7616 4048 7616 0 VGND
rlabel metal1 4048 7072 4048 7072 0 VPWR
rlabel via3 6141 5644 6141 5644 0 CLK
rlabel metal3 1188 6868 1188 6868 0 D0
rlabel metal3 751 4964 751 4964 0 D1
rlabel metal3 751 3060 751 3060 0 D2
rlabel metal3 1188 1156 1188 1156 0 D3
rlabel metal2 1426 8143 1426 8143 0 EOC
rlabel metal2 4002 1588 4002 1588 0 GND
rlabel metal2 2070 8483 2070 8483 0 NRST
rlabel metal1 6808 5202 6808 5202 0 Vcomp
rlabel metal1 4508 2618 4508 2618 0 clknet_0_CLK
rlabel metal2 1610 3060 1610 3060 0 clknet_1_0__leaf_CLK
rlabel metal1 6026 5746 6026 5746 0 clknet_1_1__leaf_CLK
rlabel metal2 3910 4182 3910 4182 0 net1
rlabel metal1 3864 5882 3864 5882 0 net10
rlabel metal1 3680 2618 3680 2618 0 net16
rlabel metal1 3772 3434 3772 3434 0 net17
rlabel metal1 4416 4114 4416 4114 0 net18
rlabel metal1 4646 4182 4646 4182 0 net19
rlabel metal1 2530 3570 2530 3570 0 net2
rlabel metal1 2392 4250 2392 4250 0 net20
rlabel metal1 4462 2890 4462 2890 0 net21
rlabel metal1 1886 2992 1886 2992 0 net22
rlabel via1 4117 5882 4117 5882 0 net23
rlabel metal1 4439 5746 4439 5746 0 net3
rlabel metal1 3197 3638 3197 3638 0 net4
rlabel metal2 5474 5644 5474 5644 0 net5
rlabel metal1 3779 3094 3779 3094 0 net6
rlabel metal1 4133 4522 4133 4522 0 net7
rlabel metal1 3496 3502 3496 3502 0 net8
rlabel metal1 3818 5610 3818 5610 0 net9
<< properties >>
string FIXED_BBOX 0 0 8127 10271
<< end >>
