** sch_path: /home/ttuser/Desktop/DAC_driver.sch
.subckt DAC_driver VPWR Dn_d Dn VGND
*.PININFO Dn_d:O Dn:I VPWR:I VGND:I
XM19 Dn_d net1 VGND VGND sky130_fd_pr__nfet_01v8_lvt L=0.5 W=6 nf=3 m=1
XM20 Dn_d net1 VPWR VPWR sky130_fd_pr__pfet_01v8_lvt L=0.5 W=10 nf=5 m=1
XM27 net1 Dn VGND VGND sky130_fd_pr__nfet_01v8_lvt L=1 W=2 nf=1 m=1
XM28 net1 Dn VPWR VPWR sky130_fd_pr__pfet_01v8_lvt L=1 W=2 nf=1 m=1
.ends
.end
