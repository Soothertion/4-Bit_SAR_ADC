* NGSPICE file created from PComp.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_lvt_5W6L9D a_400_n400# a_n458_n400# a_n400_n488# a_n560_n574#
X0 a_400_n400# a_n400_n488# a_n458_n400# a_n560_n574# sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=4
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_GWB8VV a_n258_n400# w_n396_n619# a_n200_n497#
+ a_200_n400#
X0 a_200_n400# a_n200_n497# a_n258_n400# w_n396_n619# sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_YYMWFH a_n29_n400# a_n429_n497# a_429_n400# a_29_n497#
+ w_n625_n619# a_n487_n400#
X0 a_n29_n400# a_n429_n497# a_n487_n400# w_n625_n619# sky130_fd_pr__pfet_01v8_lvt ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=2
X1 a_429_n400# a_29_n497# a_n29_n400# w_n625_n619# sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=2
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_FMZK9W a_400_n200# a_n458_n200# a_n400_n288# a_n560_n374#
X0 a_400_n200# a_n400_n288# a_n458_n200# a_n560_n374# sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=4
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_TZF6Y6 w_n246_n269# a_n108_n50# a_50_n50# a_n50_n147#
X0 a_50_n50# a_n50_n147# a_n108_n50# w_n246_n269# sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_SBHCTW a_50_n61# a_n50_n149# a_n210_n235# a_n108_n61#
X0 a_50_n61# a_n50_n149# a_n108_n61# a_n210_n235# sky130_fd_pr__nfet_01v8_lvt ad=0.1769 pd=1.8 as=0.1769 ps=1.8 w=0.61 l=0.5
.ends

.subckt PComp VPWR Vref Vin Vcomp_p VGND
XXM1 netml VGND netml VGND sky130_fd_pr__nfet_01v8_lvt_5W6L9D
XXM2 netml2 VPWR Vref VPWR sky130_fd_pr__pfet_01v8_lvt_GWB8VV
XXM3 VGND netml2 netml2 VGND sky130_fd_pr__nfet_01v8_lvt_5W6L9D
XXM4 n1 n1 VPWR n1 VPWR VPWR sky130_fd_pr__pfet_01v8_lvt_YYMWFH
XXM6 VGND m1_6268_n296# netml VGND sky130_fd_pr__nfet_01v8_lvt_FMZK9W
XXM7 VGND n1 netml2 VGND sky130_fd_pr__nfet_01v8_lvt_FMZK9W
XXM8 VPWR Vcomp_p VPWR m1_6268_n296# sky130_fd_pr__pfet_01v8_lvt_TZF6Y6
XXM9 VPWR VPWR Vin netml sky130_fd_pr__pfet_01v8_lvt_GWB8VV
Xsky130_fd_pr__pfet_01v8_lvt_YYMWFH_0 m1_6268_n296# n1 VPWR n1 VPWR VPWR sky130_fd_pr__pfet_01v8_lvt_YYMWFH
XXM10 Vcomp_p m1_6268_n296# VGND VGND sky130_fd_pr__nfet_01v8_lvt_SBHCTW
.ends

