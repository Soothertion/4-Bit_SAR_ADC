magic
tech sky130A
magscale 1 2
timestamp 1739891334
<< nwell >>
rect -562 -419 562 419
<< pmoslvt >>
rect -366 -200 -266 200
rect -208 -200 -108 200
rect -50 -200 50 200
rect 108 -200 208 200
rect 266 -200 366 200
<< pdiff >>
rect -424 188 -366 200
rect -424 -188 -412 188
rect -378 -188 -366 188
rect -424 -200 -366 -188
rect -266 188 -208 200
rect -266 -188 -254 188
rect -220 -188 -208 188
rect -266 -200 -208 -188
rect -108 188 -50 200
rect -108 -188 -96 188
rect -62 -188 -50 188
rect -108 -200 -50 -188
rect 50 188 108 200
rect 50 -188 62 188
rect 96 -188 108 188
rect 50 -200 108 -188
rect 208 188 266 200
rect 208 -188 220 188
rect 254 -188 266 188
rect 208 -200 266 -188
rect 366 188 424 200
rect 366 -188 378 188
rect 412 -188 424 188
rect 366 -200 424 -188
<< pdiffc >>
rect -412 -188 -378 188
rect -254 -188 -220 188
rect -96 -188 -62 188
rect 62 -188 96 188
rect 220 -188 254 188
rect 378 -188 412 188
<< nsubdiff >>
rect -526 349 -430 383
rect 430 349 526 383
rect -526 287 -492 349
rect 492 287 526 349
rect -526 -349 -492 -287
rect 492 -349 526 -287
rect -526 -383 -430 -349
rect 430 -383 526 -349
<< nsubdiffcont >>
rect -430 349 430 383
rect -526 -287 -492 287
rect 492 -287 526 287
rect -430 -383 430 -349
<< poly >>
rect -366 281 -266 297
rect -366 247 -350 281
rect -282 247 -266 281
rect -366 200 -266 247
rect -208 281 -108 297
rect -208 247 -192 281
rect -124 247 -108 281
rect -208 200 -108 247
rect -50 281 50 297
rect -50 247 -34 281
rect 34 247 50 281
rect -50 200 50 247
rect 108 281 208 297
rect 108 247 124 281
rect 192 247 208 281
rect 108 200 208 247
rect 266 281 366 297
rect 266 247 282 281
rect 350 247 366 281
rect 266 200 366 247
rect -366 -247 -266 -200
rect -366 -281 -350 -247
rect -282 -281 -266 -247
rect -366 -297 -266 -281
rect -208 -247 -108 -200
rect -208 -281 -192 -247
rect -124 -281 -108 -247
rect -208 -297 -108 -281
rect -50 -247 50 -200
rect -50 -281 -34 -247
rect 34 -281 50 -247
rect -50 -297 50 -281
rect 108 -247 208 -200
rect 108 -281 124 -247
rect 192 -281 208 -247
rect 108 -297 208 -281
rect 266 -247 366 -200
rect 266 -281 282 -247
rect 350 -281 366 -247
rect 266 -297 366 -281
<< polycont >>
rect -350 247 -282 281
rect -192 247 -124 281
rect -34 247 34 281
rect 124 247 192 281
rect 282 247 350 281
rect -350 -281 -282 -247
rect -192 -281 -124 -247
rect -34 -281 34 -247
rect 124 -281 192 -247
rect 282 -281 350 -247
<< locali >>
rect -526 349 -430 383
rect 430 349 526 383
rect -526 287 -492 349
rect 492 287 526 349
rect -366 247 -350 281
rect -282 247 -266 281
rect -208 247 -192 281
rect -124 247 -108 281
rect -50 247 -34 281
rect 34 247 50 281
rect 108 247 124 281
rect 192 247 208 281
rect 266 247 282 281
rect 350 247 366 281
rect -412 188 -378 204
rect -412 -204 -378 -188
rect -254 188 -220 204
rect -254 -204 -220 -188
rect -96 188 -62 204
rect -96 -204 -62 -188
rect 62 188 96 204
rect 62 -204 96 -188
rect 220 188 254 204
rect 220 -204 254 -188
rect 378 188 412 204
rect 378 -204 412 -188
rect -366 -281 -350 -247
rect -282 -281 -266 -247
rect -208 -281 -192 -247
rect -124 -281 -108 -247
rect -50 -281 -34 -247
rect 34 -281 50 -247
rect 108 -281 124 -247
rect 192 -281 208 -247
rect 266 -281 282 -247
rect 350 -281 366 -247
rect -526 -349 -492 -287
rect 492 -349 526 -287
rect -526 -383 -430 -349
rect 430 -383 526 -349
<< viali >>
rect -350 247 -282 281
rect -192 247 -124 281
rect -34 247 34 281
rect 124 247 192 281
rect 282 247 350 281
rect -412 -188 -378 188
rect -254 -188 -220 188
rect -96 -188 -62 188
rect 62 -188 96 188
rect 220 -188 254 188
rect 378 -188 412 188
rect -350 -281 -282 -247
rect -192 -281 -124 -247
rect -34 -281 34 -247
rect 124 -281 192 -247
rect 282 -281 350 -247
<< metal1 >>
rect -362 281 -270 287
rect -362 247 -350 281
rect -282 247 -270 281
rect -362 241 -270 247
rect -204 281 -112 287
rect -204 247 -192 281
rect -124 247 -112 281
rect -204 241 -112 247
rect -46 281 46 287
rect -46 247 -34 281
rect 34 247 46 281
rect -46 241 46 247
rect 112 281 204 287
rect 112 247 124 281
rect 192 247 204 281
rect 112 241 204 247
rect 270 281 362 287
rect 270 247 282 281
rect 350 247 362 281
rect 270 241 362 247
rect -418 188 -372 200
rect -418 -188 -412 188
rect -378 -188 -372 188
rect -418 -200 -372 -188
rect -260 188 -214 200
rect -260 -188 -254 188
rect -220 -188 -214 188
rect -260 -200 -214 -188
rect -102 188 -56 200
rect -102 -188 -96 188
rect -62 -188 -56 188
rect -102 -200 -56 -188
rect 56 188 102 200
rect 56 -188 62 188
rect 96 -188 102 188
rect 56 -200 102 -188
rect 214 188 260 200
rect 214 -188 220 188
rect 254 -188 260 188
rect 214 -200 260 -188
rect 372 188 418 200
rect 372 -188 378 188
rect 412 -188 418 188
rect 372 -200 418 -188
rect -362 -247 -270 -241
rect -362 -281 -350 -247
rect -282 -281 -270 -247
rect -362 -287 -270 -281
rect -204 -247 -112 -241
rect -204 -281 -192 -247
rect -124 -281 -112 -247
rect -204 -287 -112 -281
rect -46 -247 46 -241
rect -46 -281 -34 -247
rect 34 -281 46 -247
rect -46 -287 46 -281
rect 112 -247 204 -241
rect 112 -281 124 -247
rect 192 -281 204 -247
rect 112 -287 204 -281
rect 270 -247 362 -241
rect 270 -281 282 -247
rect 350 -281 362 -247
rect 270 -287 362 -281
<< properties >>
string FIXED_BBOX -509 -366 509 366
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 2.0 l 0.5 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
