magic
tech sky130A
magscale 1 2
timestamp 1739974557
<< locali >>
rect 7788 1866 8201 1868
rect 2398 1797 8201 1866
rect 2398 1699 2457 1797
rect 8152 1699 8201 1797
rect 2398 1566 8201 1699
rect 2398 399 2826 1566
rect 4158 399 4639 1566
rect 6883 1066 8200 1566
rect 6884 680 7387 1066
rect 7733 680 8200 1066
rect 6884 400 8200 680
rect 6884 399 7387 400
rect 2507 398 2741 399
rect 2402 -1227 2835 -76
rect 4959 -1227 5416 -80
rect 6796 -88 7395 -84
rect 6796 -440 8203 -88
rect 6796 -809 7395 -440
rect 7737 -809 8200 -440
rect 6796 -1227 8200 -809
rect 2401 -1354 8201 -1227
rect 2401 -1452 2473 -1354
rect 8168 -1452 8201 -1354
rect 2401 -1502 8201 -1452
<< viali >>
rect 2457 1699 8152 1797
rect 2473 -1452 8168 -1354
<< metal1 >>
rect 2398 1797 8198 1866
rect 2398 1699 2457 1797
rect 8152 1699 8198 1797
rect 2398 1668 8198 1699
rect 2398 1599 4299 1668
rect 4528 1654 8198 1668
rect 4528 1600 7008 1654
rect 7186 1600 8198 1654
rect 4528 1599 8198 1600
rect 2398 1581 8198 1599
rect 2481 1574 2696 1581
rect 3095 1499 3227 1504
rect 2961 1445 2971 1499
rect 3332 1445 3342 1499
rect 2872 668 2882 900
rect 2938 668 2948 900
rect 3095 546 3227 1445
rect 3376 1314 3602 1581
rect 3651 1447 3661 1501
rect 4022 1447 4032 1501
rect 3364 1153 3622 1314
rect 3364 908 3624 1153
rect 3365 862 3624 908
rect 3769 541 3901 1447
rect 4872 1363 5068 1503
rect 4051 912 4500 1210
rect 4872 1192 4966 1363
rect 5026 1192 5068 1363
rect 4704 944 4714 1122
rect 4768 944 4778 1122
rect 4237 320 4499 912
rect 4872 544 5068 1192
rect 5337 1363 5525 1503
rect 5337 1193 5378 1363
rect 5448 1193 5525 1363
rect 5163 643 5173 867
rect 5226 643 5236 867
rect 5337 861 5525 1193
rect 6004 1362 6195 1501
rect 6004 1189 6050 1362
rect 6109 1189 6195 1362
rect 5592 943 5602 1124
rect 5664 943 5674 1124
rect 5848 937 5858 1121
rect 5912 937 5922 1121
rect 5337 669 5374 861
rect 5452 669 5525 861
rect 5337 546 5525 669
rect 6004 547 6195 1189
rect 6465 1360 6656 1503
rect 6465 1189 6544 1360
rect 6596 1189 6656 1360
rect 6307 639 6317 851
rect 6376 639 6386 851
rect 6465 549 6656 1189
rect 6742 937 6752 1122
rect 6805 937 6815 1122
rect 7138 910 7277 1581
rect 7138 832 7498 910
rect 7534 753 7582 1000
rect 7624 889 8122 908
rect 7624 835 7881 889
rect 8107 835 8122 889
rect 7624 830 8122 835
rect 4237 159 7127 320
rect 7534 281 7586 753
rect 4242 148 7127 159
rect 5042 147 7127 148
rect 2862 -673 2872 -450
rect 2932 -673 2942 -450
rect 3198 -467 3502 -227
rect 3198 -658 3243 -467
rect 3330 -658 3502 -467
rect 3198 -1164 3502 -658
rect 4302 -549 4606 -223
rect 4302 -553 4865 -549
rect 5042 -553 5243 147
rect 5553 -294 5563 -233
rect 5931 -294 5941 -233
rect 6268 -296 6278 -233
rect 6649 -296 6659 -233
rect 3767 -1092 4022 -837
rect 4302 -860 5247 -553
rect 5438 -814 5448 -551
rect 5504 -601 5514 -551
rect 5504 -800 6016 -601
rect 6189 -797 6693 -599
rect 6899 -603 7127 147
rect 7326 273 7586 281
rect 7326 109 7369 273
rect 7446 109 7586 273
rect 7326 93 7586 109
rect 7534 -528 7586 93
rect 7535 -543 7586 -528
rect 6699 -797 7127 -603
rect 7163 -679 7502 -584
rect 6189 -799 7127 -797
rect 5504 -814 5514 -800
rect 4302 -872 4865 -860
rect 2500 -1257 2736 -1242
rect 3818 -1257 3975 -1092
rect 4302 -1160 4606 -872
rect 5563 -1257 5935 -1123
rect 6276 -1257 6645 -1122
rect 7166 -1257 7317 -679
rect 7540 -722 7586 -543
rect 7629 -599 8119 -589
rect 7629 -675 7889 -599
rect 8099 -675 8119 -599
rect 7629 -682 8119 -675
rect 7535 -764 7586 -722
rect 2402 -1354 8198 -1257
rect 2402 -1452 2473 -1354
rect 8168 -1452 8198 -1354
rect 2402 -1500 8198 -1452
<< via1 >>
rect 4299 1599 4528 1668
rect 7008 1600 7186 1654
rect 2971 1445 3332 1499
rect 2882 668 2938 900
rect 3661 1447 4022 1501
rect 4966 1192 5026 1363
rect 4714 944 4768 1122
rect 5378 1193 5448 1363
rect 5173 643 5226 867
rect 6050 1189 6109 1362
rect 5602 943 5664 1124
rect 5858 937 5912 1121
rect 5374 669 5452 861
rect 6544 1189 6596 1360
rect 6317 639 6376 851
rect 6752 937 6805 1122
rect 7881 835 8107 889
rect 2872 -673 2932 -450
rect 3243 -658 3330 -467
rect 5563 -294 5931 -233
rect 6278 -296 6649 -233
rect 5448 -814 5504 -551
rect 7369 109 7446 273
rect 7889 -675 8099 -599
<< metal2 >>
rect 3001 1509 3294 2236
rect 3691 1511 3984 2241
rect 4299 1675 4528 1678
rect 4293 1668 4542 1675
rect 4293 1599 4299 1668
rect 4528 1599 4542 1668
rect 7008 1662 7186 1664
rect 2971 1499 3332 1509
rect 2971 1435 3332 1445
rect 3661 1501 4022 1511
rect 3661 1437 4022 1447
rect 4293 1121 4542 1599
rect 6996 1654 7200 1662
rect 6996 1600 7008 1654
rect 7186 1600 7200 1654
rect 4948 1375 5460 1377
rect 4948 1363 6626 1375
rect 4948 1192 4966 1363
rect 5026 1193 5378 1363
rect 5448 1362 6626 1363
rect 5448 1193 6050 1362
rect 5026 1192 6050 1193
rect 4948 1189 6050 1192
rect 6109 1360 6626 1362
rect 6109 1189 6544 1360
rect 6596 1189 6626 1360
rect 4948 1183 6626 1189
rect 4966 1182 5026 1183
rect 5378 1182 6626 1183
rect 6035 1180 6626 1182
rect 6050 1179 6109 1180
rect 6544 1179 6596 1180
rect 4714 1126 4768 1132
rect 5602 1126 5664 1134
rect 4714 1124 5668 1126
rect 5858 1124 5912 1131
rect 6752 1124 6805 1132
rect 4714 1122 5602 1124
rect 4293 944 4714 1121
rect 4768 944 5602 1122
rect 4293 943 4542 944
rect 4714 943 5602 944
rect 5664 943 5668 1124
rect 4714 941 5668 943
rect 5857 1122 6808 1124
rect 6996 1122 7200 1600
rect 5857 1121 6752 1122
rect 4714 934 4768 941
rect 5602 933 5664 941
rect 5857 937 5858 1121
rect 5912 937 6752 1121
rect 6805 937 7200 1122
rect 5857 934 7200 937
rect 5857 933 6808 934
rect 5858 927 5912 933
rect 6752 927 6805 933
rect 2882 900 2938 910
rect 2547 899 2882 900
rect 2505 739 2882 899
rect 2506 668 2882 739
rect 2938 668 2939 900
rect 7881 894 8107 899
rect 7881 889 8115 894
rect 5173 874 5226 877
rect 5510 874 5553 875
rect 2506 663 2939 668
rect 5171 867 5553 874
rect 2506 372 2742 663
rect 2882 658 2938 663
rect 5171 643 5173 867
rect 5226 861 5553 867
rect 5226 669 5374 861
rect 5452 720 5553 861
rect 6317 854 6376 861
rect 6317 851 6651 854
rect 5452 669 5555 720
rect 5226 643 5555 669
rect 5171 637 5555 643
rect 5173 633 5226 637
rect 2504 354 2742 372
rect 2502 220 2742 354
rect 5337 499 5555 637
rect 6376 639 6651 851
rect 6317 636 6651 639
rect 6317 629 6376 636
rect 5337 332 5797 499
rect 5537 331 5797 332
rect 2506 197 2742 220
rect 5002 197 5376 198
rect 2506 64 5376 197
rect 2506 4 5380 64
rect 2506 -59 2742 4
rect 2507 -443 2741 -59
rect 2872 -443 2932 -440
rect 2506 -447 2939 -443
rect 2506 -450 3356 -447
rect 2506 -673 2872 -450
rect 2932 -467 3356 -450
rect 2932 -658 3243 -467
rect 3330 -658 3356 -467
rect 2932 -673 3356 -658
rect 2506 -680 3356 -673
rect 2851 -683 3356 -680
rect 5188 -549 5380 4
rect 5561 -101 5797 331
rect 6430 287 6651 636
rect 8107 835 8115 889
rect 6430 273 7462 287
rect 6430 109 7369 273
rect 7446 109 7462 273
rect 6430 90 7462 109
rect 6430 -30 6651 90
rect 5561 -233 5934 -101
rect 5561 -294 5563 -233
rect 5931 -294 5934 -233
rect 5561 -296 5934 -294
rect 6274 -233 6651 -30
rect 6274 -296 6278 -233
rect 6649 -296 6651 -233
rect 5563 -304 5931 -296
rect 6274 -300 6651 -296
rect 6278 -306 6649 -300
rect 5448 -549 5504 -541
rect 5188 -551 5508 -549
rect 5188 -814 5448 -551
rect 5504 -814 5508 -551
rect 7881 -599 8115 835
rect 7881 -675 7889 -599
rect 8099 -675 8115 -599
rect 7881 -679 8115 -675
rect 7889 -685 8099 -679
rect 5188 -816 5508 -814
rect 5290 -817 5508 -816
rect 5448 -824 5504 -817
use sky130_fd_pr__pfet_01v8_lvt_YYMWFH  sky130_fd_pr__pfet_01v8_lvt_YYMWFH_0
timestamp 1739974041
transform 1 0 6334 0 1 1020
box -625 -619 625 619
use sky130_fd_pr__nfet_01v8_lvt_5W6L9D  XM1
timestamp 1739436521
transform 1 0 4437 0 1 -691
box -596 -610 596 610
use sky130_fd_pr__pfet_01v8_lvt_GWB8VV  XM2
timestamp 1739902357
transform 1 0 3152 0 1 1019
box -396 -619 396 619
use sky130_fd_pr__nfet_01v8_lvt_5W6L9D  XM3
timestamp 1739436521
transform 1 0 3351 0 1 -691
box -596 -610 596 610
use sky130_fd_pr__pfet_01v8_lvt_YYMWFH  XM4
timestamp 1739974041
transform 1 0 5190 0 1 1020
box -625 -619 625 619
use sky130_fd_pr__nfet_01v8_lvt_FMZK9W  XM6
timestamp 1739902357
transform 0 1 6461 -1 0 -710
box -596 -410 596 410
use sky130_fd_pr__nfet_01v8_lvt_FMZK9W  XM7
timestamp 1739902357
transform 0 1 5747 -1 0 -710
box -596 -410 596 410
use sky130_fd_pr__pfet_01v8_lvt_TZF6Y6  XM8
timestamp 1739902357
transform -1 0 7560 0 1 871
box -246 -269 246 269
use sky130_fd_pr__pfet_01v8_lvt_GWB8VV  XM9
timestamp 1739902357
transform 1 0 3838 0 1 1019
box -396 -619 396 619
use sky130_fd_pr__nfet_01v8_lvt_SBHCTW  XM10
timestamp 1739436521
transform 1 0 7565 0 1 -633
box -246 -271 246 271
<< labels >>
flabel metal1 2585 -1480 2785 -1280 0 FreeSans 256 0 0 0 VGND
port 4 nsew
flabel metal1 2465 1628 2665 1828 0 FreeSans 256 0 0 0 VPWR
port 0 nsew
flabel metal2 3036 2008 3236 2208 0 FreeSans 256 0 0 0 Vref
port 1 nsew
flabel metal2 3739 1995 3939 2195 0 FreeSans 256 0 0 0 Vin
port 2 nsew
flabel metal2 7892 -2 8092 198 0 FreeSans 256 0 0 0 Vcomp_p
port 3 nsew
flabel metal2 2540 16 3056 174 0 FreeSans 800 0 0 0 netml2
flabel metal1 4252 226 4450 338 0 FreeSans 640 0 0 0 netml
flabel metal2 5578 -15 5786 143 0 FreeSans 800 0 0 0 n1
<< end >>
