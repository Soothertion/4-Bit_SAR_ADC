magic
tech sky130A
timestamp 1739797948
<< pwell >>
rect -148 -305 148 305
<< nmoslvt >>
rect -50 -200 50 200
<< ndiff >>
rect -79 194 -50 200
rect -79 -194 -73 194
rect -56 -194 -50 194
rect -79 -200 -50 -194
rect 50 194 79 200
rect 50 -194 56 194
rect 73 -194 79 194
rect 50 -200 79 -194
<< ndiffc >>
rect -73 -194 -56 194
rect 56 -194 73 194
<< psubdiff >>
rect -130 270 -82 287
rect 82 270 130 287
rect -130 239 -113 270
rect 113 239 130 270
rect -130 -270 -113 -239
rect 113 -270 130 -239
rect -130 -287 -82 -270
rect 82 -287 130 -270
<< psubdiffcont >>
rect -82 270 82 287
rect -130 -239 -113 239
rect 113 -239 130 239
rect -82 -287 82 -270
<< poly >>
rect -50 236 50 244
rect -50 219 -42 236
rect 42 219 50 236
rect -50 200 50 219
rect -50 -219 50 -200
rect -50 -236 -42 -219
rect 42 -236 50 -219
rect -50 -244 50 -236
<< polycont >>
rect -42 219 42 236
rect -42 -236 42 -219
<< locali >>
rect -130 270 -82 287
rect 82 270 130 287
rect -130 239 -113 270
rect 113 239 130 270
rect -50 219 -42 236
rect 42 219 50 236
rect -73 194 -56 202
rect -73 -202 -56 -194
rect 56 194 73 202
rect 56 -202 73 -194
rect -50 -236 -42 -219
rect 42 -236 50 -219
rect -130 -270 -113 -239
rect 113 -270 130 -239
rect -130 -287 -82 -270
rect 82 -287 130 -270
<< viali >>
rect -42 219 42 236
rect -73 -194 -56 194
rect 56 -194 73 194
rect -42 -236 42 -219
<< metal1 >>
rect -48 236 48 239
rect -48 219 -42 236
rect 42 219 48 236
rect -48 216 48 219
rect -76 194 -53 200
rect -76 -194 -73 194
rect -56 -194 -53 194
rect -76 -200 -53 -194
rect 53 194 76 200
rect 53 -194 56 194
rect 73 -194 76 194
rect 53 -200 76 -194
rect -48 -219 48 -216
rect -48 -236 -42 -219
rect 42 -236 48 -219
rect -48 -239 48 -236
<< properties >>
string FIXED_BBOX -121 -278 121 278
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 4.0 l 1.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
