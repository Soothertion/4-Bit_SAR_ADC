magic
tech sky130A
magscale 1 2
timestamp 1739891334
<< locali >>
rect 760 1145 2458 1185
rect 760 984 1006 1145
rect 2407 984 2458 1145
rect 760 873 2458 984
rect 760 141 881 873
rect 2349 141 2458 873
rect 760 -870 882 -156
rect 2032 -870 2123 -157
rect 760 -942 2123 -870
rect 759 -986 2123 -942
rect 759 -1140 1007 -986
rect 2072 -1140 2123 -986
rect 759 -1182 2123 -1140
<< viali >>
rect 1006 984 2407 1145
rect 1007 -1140 2072 -986
<< metal1 >>
rect 782 1145 2437 1164
rect 782 1088 1006 1145
rect 782 964 899 1088
rect 889 954 899 964
rect 952 984 1006 1088
rect 2407 984 2437 1145
rect 952 968 1385 984
rect 1437 971 1753 984
rect 1805 971 2069 984
rect 2121 971 2437 984
rect 1437 968 2437 971
rect 952 964 2437 968
rect 952 954 962 964
rect 929 340 939 710
rect 991 340 1001 710
rect 1076 87 1136 807
rect 1514 739 1570 807
rect 1672 739 1728 807
rect 1830 739 1886 807
rect 1988 739 2044 807
rect 2146 739 2202 807
rect 1217 336 1326 714
rect 1413 340 1423 709
rect 1475 340 1485 709
rect 1286 89 1326 336
rect 1514 312 1556 739
rect 1585 341 1595 710
rect 1647 341 1657 710
rect 1686 312 1714 739
rect 1743 343 1753 713
rect 1805 343 1815 713
rect 1844 312 1872 739
rect 1901 343 1911 708
rect 1963 343 1973 708
rect 2002 312 2030 739
rect 2059 340 2069 710
rect 2121 340 2131 710
rect 2160 312 2188 739
rect 2217 341 2227 708
rect 2279 341 2289 708
rect 1514 89 1570 312
rect 1672 89 1728 312
rect 1830 197 1886 312
rect 1988 197 2044 312
rect 2146 197 2202 312
rect 1830 145 2202 197
rect 1830 89 1886 145
rect 1070 -105 1080 87
rect 1132 -105 1142 87
rect 1286 9 1886 89
rect 930 -717 940 -346
rect 992 -717 1002 -346
rect 1076 -805 1136 -105
rect 1286 -343 1326 9
rect 1217 -721 1326 -343
rect 1514 -318 1570 9
rect 1672 -318 1728 9
rect 1830 -318 1886 9
rect 1414 -717 1424 -347
rect 1476 -717 1486 -347
rect 1514 -746 1556 -318
rect 1585 -717 1595 -347
rect 1647 -717 1657 -347
rect 1686 -746 1714 -318
rect 1743 -716 1753 -347
rect 1805 -716 1815 -347
rect 1844 -745 1872 -318
rect 1901 -716 1911 -347
rect 1963 -716 1973 -347
rect 1844 -746 1886 -745
rect 1514 -805 1570 -746
rect 1672 -805 1728 -746
rect 1830 -805 1886 -746
rect 785 -965 2089 -962
rect 785 -967 1385 -965
rect 785 -1079 899 -967
rect 951 -986 1385 -967
rect 1437 -967 2089 -965
rect 1437 -986 1752 -967
rect 1804 -986 2089 -967
rect 951 -1079 1007 -986
rect 785 -1140 1007 -1079
rect 2072 -1140 2089 -986
rect 785 -1162 2089 -1140
<< via1 >>
rect 899 954 952 1088
rect 1385 984 1437 1075
rect 1753 984 1805 1077
rect 2069 984 2121 1077
rect 1385 968 1437 984
rect 1753 971 1805 984
rect 2069 971 2121 984
rect 939 340 991 710
rect 1423 340 1475 709
rect 1595 341 1647 710
rect 1753 343 1805 713
rect 1911 343 1963 708
rect 2069 340 2121 710
rect 2227 341 2279 708
rect 1080 -105 1132 87
rect 940 -717 992 -346
rect 1424 -717 1476 -347
rect 1595 -717 1647 -347
rect 1753 -716 1805 -347
rect 1911 -716 1963 -347
rect 899 -1079 951 -967
rect 1385 -986 1437 -965
rect 1752 -986 1804 -967
rect 1385 -1076 1437 -986
rect 1752 -1079 1804 -986
<< metal2 >>
rect 899 1091 952 1098
rect 895 1088 955 1091
rect 895 954 899 1088
rect 952 954 955 1088
rect 1385 1078 1437 1085
rect 895 720 955 954
rect 1381 1075 1441 1078
rect 1381 968 1385 1075
rect 1437 968 1441 1075
rect 895 714 991 720
rect 1381 719 1441 968
rect 1753 1077 1805 1087
rect 1381 714 1475 719
rect 895 710 995 714
rect 895 340 939 710
rect 991 340 995 710
rect 895 336 995 340
rect 1381 709 1481 714
rect 1381 340 1423 709
rect 1475 340 1481 709
rect 1381 336 1481 340
rect 1595 710 1647 720
rect 939 330 991 336
rect 1423 330 1475 336
rect 1080 92 1132 97
rect 936 87 1136 92
rect 936 -105 1080 87
rect 1132 -105 1136 87
rect 1595 -23 1647 341
rect 1753 713 1805 971
rect 2069 1077 2121 1087
rect 1753 333 1805 343
rect 1911 708 1963 718
rect 1911 -23 1963 343
rect 2069 710 2121 971
rect 2069 330 2121 340
rect 2227 708 2279 718
rect 2227 96 2279 341
rect 2227 -23 2427 96
rect 1594 -103 2427 -23
rect 936 -108 1136 -105
rect 1080 -115 1132 -108
rect 940 -343 992 -336
rect 1424 -343 1476 -337
rect 895 -346 995 -343
rect 895 -717 940 -346
rect 992 -717 995 -346
rect 895 -721 995 -717
rect 1381 -347 1481 -343
rect 1381 -717 1424 -347
rect 1476 -717 1481 -347
rect 1381 -721 1481 -717
rect 1595 -347 1647 -103
rect 895 -727 992 -721
rect 1381 -727 1476 -721
rect 895 -967 955 -727
rect 895 -1079 899 -967
rect 951 -1079 955 -967
rect 895 -1085 955 -1079
rect 1381 -965 1441 -727
rect 1595 -739 1647 -717
rect 1753 -347 1805 -337
rect 1753 -957 1805 -716
rect 1911 -347 1963 -103
rect 2227 -104 2427 -103
rect 1911 -726 1963 -716
rect 1381 -1076 1385 -965
rect 1437 -1076 1441 -965
rect 1381 -1081 1441 -1076
rect 1752 -967 1805 -957
rect 1804 -1079 1805 -967
rect 899 -1089 951 -1085
rect 1385 -1086 1437 -1081
rect 1752 -1089 1804 -1079
use sky130_fd_pr__nfet_01v8_lvt_56BWKP  XM19
timestamp 1739891334
transform 1 0 1700 0 1 -532
box -404 -410 404 410
use sky130_fd_pr__pfet_01v8_lvt_X33VY6  XM20
timestamp 1739891334
transform 1 0 1858 0 1 525
box -562 -419 562 419
use sky130_fd_pr__nfet_01v8_lvt_QGMAL3  XM27
timestamp 1739891334
transform 1 0 1106 0 1 -532
box -296 -410 296 410
use sky130_fd_pr__pfet_01v8_lvt_3VC8VM  XM28
timestamp 1739891334
transform 1 0 1106 0 1 525
box -296 -419 296 419
<< labels >>
flabel metal1 785 -1162 985 -962 0 FreeSans 256 0 0 0 VGND
port 3 nsew
flabel metal1 782 964 982 1164 0 FreeSans 256 0 0 0 VPWR
port 2 nsew
flabel metal2 936 -108 1136 92 0 FreeSans 256 0 0 0 Dn
port 1 nsew
flabel metal2 2227 -104 2427 96 0 FreeSans 256 0 0 0 Dn_d
port 0 nsew
<< end >>
