magic
tech sky130A
magscale 1 2
timestamp 1739900237
<< pwell >>
rect -201 -1782 201 1782
<< psubdiff >>
rect -165 1712 -69 1746
rect 69 1712 165 1746
rect -165 1650 -131 1712
rect 131 1650 165 1712
rect -165 -1712 -131 -1650
rect 131 -1712 165 -1650
rect -165 -1746 -69 -1712
rect 69 -1746 165 -1712
<< psubdiffcont >>
rect -69 1712 69 1746
rect -165 -1650 -131 1650
rect 131 -1650 165 1650
rect -69 -1746 69 -1712
<< xpolycontact >>
rect -35 1184 35 1616
rect -35 -1616 35 -1184
<< ppolyres >>
rect -35 -1184 35 1184
<< locali >>
rect -165 1712 -69 1746
rect 69 1712 165 1746
rect -165 1650 -131 1712
rect 131 1650 165 1712
rect -165 -1712 -131 -1650
rect 131 -1712 165 -1650
rect -165 -1746 -69 -1712
rect 69 -1746 165 -1712
<< viali >>
rect -19 1201 19 1598
rect -19 -1598 19 -1201
<< metal1 >>
rect -25 1598 25 1610
rect -25 1201 -19 1598
rect 19 1201 25 1598
rect -25 1189 25 1201
rect -25 -1201 25 -1189
rect -25 -1598 -19 -1201
rect 19 -1598 25 -1201
rect -25 -1610 25 -1598
<< properties >>
string FIXED_BBOX -148 -1729 148 1729
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 12.0 m 1 nx 1 wmin 0.350 lmin 0.50 rho 319.8 val 12.077k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
