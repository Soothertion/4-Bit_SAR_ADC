magic
tech sky130A
magscale 1 2
timestamp 1739797948
<< metal4 >>
rect -1349 2539 1349 2580
rect -1349 -2539 1093 2539
rect 1329 -2539 1349 2539
rect -1349 -2580 1349 -2539
<< via4 >>
rect 1093 -2539 1329 2539
<< mimcap2 >>
rect -1269 2460 731 2500
rect -1269 -2460 -1229 2460
rect 691 -2460 731 2460
rect -1269 -2500 731 -2460
<< mimcap2contact >>
rect -1229 -2460 691 2460
<< metal5 >>
rect 1051 2539 1371 2581
rect -1253 2460 715 2484
rect -1253 -2460 -1229 2460
rect 691 -2460 715 2460
rect -1253 -2484 715 -2460
rect 1051 -2539 1093 2539
rect 1329 -2539 1371 2539
rect 1051 -2581 1371 -2539
<< properties >>
string FIXED_BBOX -1349 -2580 811 2580
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 10.0 l 25.0 val 513.299 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
