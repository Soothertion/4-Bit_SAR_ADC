magic
tech sky130A
magscale 1 2
timestamp 1739900237
<< locali >>
rect -1445 3424 250 3537
rect -1445 3411 251 3424
rect -1445 3354 -931 3411
rect -1445 1689 -1293 3354
rect -1144 1689 -931 3354
rect -1445 1430 -931 1689
rect -673 1430 -529 3411
rect -271 1430 -127 3411
rect 132 1430 251 3411
rect -1445 1368 251 1430
rect -1445 1291 619 1368
rect -1445 1286 620 1291
rect -1445 -1621 -1332 1286
rect -1445 -2026 -1177 -1621
rect -1075 -1812 -931 1286
rect -675 -1732 -529 1286
rect -271 -1732 -127 1286
rect 132 -1702 275 1286
rect 132 -1731 273 -1702
rect 533 -1771 620 1286
rect -1445 -2076 -1332 -2026
<< viali >>
rect -1293 1689 -1144 3354
<< metal1 >>
rect -1319 3354 -1119 3373
rect -1319 1689 -1293 3354
rect -1144 1689 -1119 3354
rect -838 2902 -828 3292
rect -776 2902 -766 3292
rect -436 2902 -426 3292
rect -374 2902 -364 3292
rect -34 2902 -24 3292
rect 28 2902 38 3292
rect -1319 1466 -1119 1689
rect -838 1543 -828 1933
rect -776 1543 -766 1933
rect -436 1543 -426 1933
rect -374 1543 -364 1933
rect -34 1543 -24 1933
rect 28 1543 38 1933
rect -1237 780 -1227 1170
rect -1175 780 -1165 1170
rect -847 780 -837 1170
rect -785 780 -775 1170
rect -436 778 -426 1168
rect -374 778 -364 1168
rect -34 778 -24 1168
rect 28 778 38 1168
rect 368 778 378 1168
rect 430 778 440 1168
rect -838 -1661 -828 -1271
rect -776 -1661 -766 -1271
rect -436 -1581 -426 -1191
rect -374 -1581 -364 -1191
rect -34 -1581 -24 -1191
rect 28 -1581 38 -1191
rect 368 -1621 378 -1231
rect 430 -1621 440 -1231
<< via1 >>
rect -828 2902 -776 3292
rect -426 2902 -374 3292
rect -24 2902 28 3292
rect -828 1543 -776 1933
rect -426 1543 -374 1933
rect -24 1543 28 1933
rect -1227 780 -1175 1170
rect -837 780 -785 1170
rect -426 778 -374 1168
rect -24 778 28 1168
rect 378 778 430 1168
rect -828 -1661 -776 -1271
rect -426 -1581 -374 -1191
rect -24 -1581 28 -1191
rect 378 -1621 430 -1231
<< metal2 >>
rect -828 3292 -776 3302
rect -426 3292 -374 3302
rect -776 2902 -578 3275
rect -828 2901 -578 2902
rect -828 2892 -776 2901
rect -828 1933 -776 1943
rect -618 1925 -578 2901
rect -24 3292 28 3302
rect -374 2908 -24 3285
rect -426 2892 -374 2902
rect -426 1933 -374 1943
rect -618 1551 -426 1925
rect -828 1180 -776 1543
rect -1227 1172 -1175 1180
rect -837 1172 -776 1180
rect -1229 1170 -776 1172
rect -1229 780 -1227 1170
rect -1175 780 -837 1170
rect -785 780 -782 1170
rect -1229 778 -782 780
rect -426 1168 -374 1543
rect -219 1162 -179 2908
rect -24 2892 28 2902
rect -24 1933 28 1943
rect 28 1547 430 1747
rect -24 1533 28 1543
rect -24 1168 28 1178
rect -219 788 -24 1162
rect -1227 770 -1175 778
rect -837 770 -785 778
rect -426 768 -374 778
rect -24 768 28 778
rect 378 1168 430 1547
rect 378 768 430 778
rect -426 -1191 -374 -1181
rect -828 -1271 -776 -1261
rect -828 -1876 -776 -1661
rect -426 -1876 -374 -1581
rect -24 -1191 28 -1181
rect 378 -1231 430 -1221
rect -24 -1876 29 -1581
rect 378 -1876 430 -1621
rect -828 -2076 -628 -1876
rect -426 -2076 -226 -1876
rect -24 -2076 176 -1876
rect 378 -2076 578 -1876
use sky130_fd_pr__res_high_po_0p35_AT4384  XR1
timestamp 1739900237
transform 1 0 -1203 0 1 -424
box -201 -1782 201 1782
use sky130_fd_pr__res_high_po_0p35_Z689S7  XR2
timestamp 1739900237
transform 1 0 -400 0 1 2420
box -201 -1062 201 1062
use sky130_fd_pr__res_high_po_0p35_Z689S7  XR3
timestamp 1739900237
transform 1 0 2 0 1 2420
box -201 -1062 201 1062
use sky130_fd_pr__res_high_po_0p35_V3ZUAZ  XR4
timestamp 1739900237
transform 1 0 -802 0 1 -244
box -201 -1602 201 1602
use sky130_fd_pr__res_high_po_0p35_GHF3PF  XR5
timestamp 1739900237
transform 1 0 -400 0 1 -204
box -201 -1562 201 1562
use sky130_fd_pr__res_high_po_0p35_GHF3PF  XR6
timestamp 1739900237
transform 1 0 2 0 1 -204
box -201 -1562 201 1562
use sky130_fd_pr__res_high_po_0p35_FFK5MY  XR7
timestamp 1739900237
transform 1 0 404 0 1 -224
box -201 -1582 201 1582
use sky130_fd_pr__res_high_po_0p35_Z689S7  XR9
timestamp 1739900237
transform 1 0 -802 0 1 2420
box -201 -1062 201 1062
<< labels >>
flabel metal2 230 1547 430 1747 0 FreeSans 256 0 0 0 Vdac
port 0 nsew
flabel metal2 -426 -2076 -226 -1876 0 FreeSans 256 0 0 0 D1
port 4 nsew
flabel metal2 -24 -2076 176 -1876 0 FreeSans 256 0 0 0 D2
port 2 nsew
flabel metal2 -828 -2076 -628 -1876 0 FreeSans 256 0 0 0 D0
port 1 nsew
flabel metal2 378 -2076 578 -1876 0 FreeSans 256 0 0 0 D3
port 3 nsew
flabel metal1 -1319 1466 -1119 1666 0 FreeSans 256 0 0 0 VGND
port 5 nsew
<< end >>
