magic
tech sky130A
magscale 1 2
timestamp 1739911419
<< pwell >>
rect 4567 -2321 4728 -1961
<< locali >>
rect 126 -190 4996 -118
rect 126 -311 403 -190
rect 4098 -311 4996 -190
rect 126 -453 4996 -311
rect 126 -1584 293 -453
rect 941 -610 1682 -453
rect 827 -999 1682 -610
rect 2616 -609 3360 -453
rect 2616 -999 3474 -609
rect 4008 -1047 4996 -453
rect 4008 -1195 4611 -1047
rect 4008 -1295 4728 -1195
rect 4008 -1480 4611 -1295
rect 4008 -1584 4190 -1480
rect -299 -1971 -165 -1784
rect 4464 -1961 4613 -1785
rect -299 -2749 -53 -1971
rect 4464 -1972 4728 -1961
rect 827 -2749 1084 -2183
rect -299 -2897 -165 -2749
rect 938 -2897 1084 -2749
rect 3214 -2750 3473 -2183
rect 4353 -2321 4728 -1972
rect 4353 -2458 4613 -2321
rect 4353 -2750 5000 -2458
rect 3214 -2897 3360 -2750
rect 4465 -2897 5000 -2750
rect -299 -3068 5000 -2897
rect -299 -3210 -22 -3068
rect 4844 -3179 5000 -3068
rect 4844 -3210 5001 -3179
rect -299 -3281 5001 -3210
<< viali >>
rect 403 -311 4098 -190
rect -22 -3210 4844 -3068
<< metal1 >>
rect 162 -190 4147 -148
rect 162 -311 403 -190
rect 4098 -311 4147 -190
rect 162 -348 4147 -311
rect 351 -998 361 -616
rect 413 -998 423 -616
rect 587 -1440 647 -542
rect 1727 -1383 1737 -1002
rect 1789 -1383 1799 -1002
rect 1876 -1445 1936 -548
rect 2099 -609 2199 -348
rect 2014 -1003 2283 -609
rect 742 -1642 802 -1445
rect 1822 -1446 1936 -1445
rect 2362 -1445 2422 -549
rect 2499 -1382 2509 -999
rect 2561 -1382 2571 -999
rect 1822 -1642 1892 -1446
rect 2362 -1447 2477 -1445
rect 2405 -1641 2477 -1447
rect 3499 -1641 3559 -1445
rect 3654 -1446 3714 -548
rect 3877 -997 3887 -614
rect 3939 -997 3949 -614
rect 735 -1694 745 -1642
rect 799 -1694 809 -1642
rect 1815 -1694 1825 -1642
rect 1888 -1694 1898 -1642
rect 2398 -1693 2408 -1641
rect 2474 -1693 2484 -1641
rect 3492 -1693 3502 -1641
rect 3556 -1693 3566 -1641
rect 4758 -1651 4810 -1148
rect 4840 -1282 4850 -1208
rect 4902 -1282 4912 -1208
rect 3877 -1703 3887 -1651
rect 3939 -1703 4810 -1651
rect 351 -1780 361 -1728
rect 413 -1780 3559 -1728
rect 128 -2797 188 -1922
rect 342 -1931 361 -1879
rect 413 -1931 432 -1879
rect 3499 -1888 3559 -1780
rect 351 -2741 361 -2359
rect 413 -2741 423 -2359
rect 586 -2797 646 -1905
rect 3499 -1924 4327 -1888
rect 1577 -1998 1677 -1987
rect 2580 -1997 2680 -1985
rect 1573 -2058 1583 -1998
rect 1671 -2058 1681 -1998
rect 2578 -2057 2588 -1997
rect 2671 -2057 2681 -1997
rect 1127 -2742 1137 -2376
rect 1189 -2742 1199 -2376
rect -27 -2833 802 -2797
rect 1577 -2833 1677 -2058
rect 2017 -2749 2281 -2371
rect 353 -2838 422 -2833
rect 2099 -3039 2199 -2749
rect 2580 -2833 2680 -2057
rect 3099 -2743 3109 -2376
rect 3161 -2743 3171 -2376
rect 3654 -2798 3714 -1924
rect 3877 -2744 3887 -2361
rect 3939 -2744 3949 -2361
rect 4112 -2798 4172 -1924
rect 4758 -2359 4810 -1703
rect 4842 -2139 4852 -1975
rect 4904 -2139 4914 -1975
rect 3499 -2834 4327 -2798
rect -254 -3068 4882 -3039
rect -254 -3210 -22 -3068
rect 4844 -3210 4882 -3068
rect -254 -3239 4882 -3210
<< via1 >>
rect 361 -998 413 -616
rect 1737 -1383 1789 -1002
rect 2509 -1382 2561 -999
rect 3887 -997 3939 -614
rect 745 -1694 799 -1642
rect 1825 -1694 1888 -1642
rect 2408 -1693 2474 -1641
rect 3502 -1693 3556 -1641
rect 4850 -1282 4902 -1208
rect 3887 -1703 3939 -1651
rect 361 -1780 413 -1728
rect 361 -1931 413 -1879
rect 361 -2741 413 -2359
rect 1583 -2058 1671 -1998
rect 2588 -2057 2671 -1997
rect 1137 -2742 1189 -2376
rect 3109 -2743 3161 -2376
rect 3887 -2744 3939 -2361
rect 4852 -2139 4904 -1975
<< metal2 >>
rect 361 -616 413 -606
rect 3887 -614 3939 -604
rect 1737 -997 1789 -992
rect 2509 -995 2561 -989
rect 361 -1728 413 -998
rect 1675 -1002 1795 -997
rect 1675 -1383 1737 -1002
rect 1789 -1383 1795 -1002
rect 1675 -1388 1795 -1383
rect 2503 -999 2623 -995
rect 2503 -1382 2509 -999
rect 2561 -1382 2623 -999
rect 2503 -1388 2623 -1382
rect 1675 -1393 1789 -1388
rect 2509 -1392 2623 -1388
rect 745 -1642 799 -1632
rect 1675 -1642 1755 -1393
rect 1825 -1642 1888 -1632
rect 2408 -1641 2474 -1631
rect 2543 -1641 2623 -1392
rect 3502 -1641 3556 -1631
rect 742 -1694 745 -1642
rect 799 -1694 1825 -1642
rect 1888 -1694 1892 -1642
rect 745 -1704 799 -1694
rect 361 -1879 413 -1780
rect 361 -2359 413 -1931
rect 1095 -1722 1892 -1694
rect 2405 -1693 2408 -1641
rect 2474 -1693 3502 -1641
rect 3556 -1693 3559 -1641
rect 3887 -1651 3939 -997
rect 4850 -1206 4902 -1198
rect 4845 -1208 4945 -1206
rect 4845 -1282 4850 -1208
rect 4902 -1282 4945 -1208
rect 4845 -1284 4945 -1282
rect 4850 -1292 4945 -1284
rect 4885 -1531 4945 -1292
rect 2405 -1721 3203 -1693
rect 3502 -1703 3556 -1693
rect 1095 -2366 1155 -1722
rect 1477 -1998 1677 -1865
rect 1477 -2058 1583 -1998
rect 1671 -2058 1677 -1998
rect 1477 -2065 1677 -2058
rect 2480 -1997 2680 -1865
rect 2480 -2057 2588 -1997
rect 2671 -2057 2680 -1997
rect 2480 -2065 2680 -2057
rect 1583 -2068 1671 -2065
rect 2588 -2067 2671 -2065
rect 3143 -2366 3203 -1721
rect 1095 -2370 1189 -2366
rect 361 -2751 413 -2741
rect 1096 -2376 1196 -2370
rect 3109 -2371 3203 -2366
rect 1096 -2742 1137 -2376
rect 1189 -2742 1196 -2376
rect 1096 -2750 1196 -2742
rect 3103 -2376 3203 -2371
rect 3103 -2743 3109 -2376
rect 3161 -2743 3203 -2376
rect 3103 -2749 3203 -2743
rect 3887 -2361 3939 -1703
rect 4884 -1731 5084 -1531
rect 4885 -1965 4945 -1731
rect 4852 -1972 4945 -1965
rect 4845 -1975 4945 -1972
rect 4845 -2139 4852 -1975
rect 4904 -2139 4945 -1975
rect 4845 -2142 4945 -2139
rect 4852 -2149 4904 -2142
rect 1137 -2752 1189 -2750
rect 3109 -2753 3161 -2749
rect 3887 -2754 3939 -2744
use sky130_fd_pr__nfet_01v8_lvt_FMZK9W  XM29
timestamp 1739902357
transform 1 0 1606 0 1 -2560
box -596 -410 596 410
use sky130_fd_pr__nfet_01v8_lvt_FMZK9W  XM30
timestamp 1739902357
transform 1 0 2692 0 1 -2560
box -596 -410 596 410
use sky130_fd_pr__pfet_01v8_lvt_3VA8VM  XM31
timestamp 1739902357
transform 1 0 1906 0 1 -999
box -296 -619 296 619
use sky130_fd_pr__pfet_01v8_lvt_3VA8VM  XM32
timestamp 1739902357
transform 1 0 2392 0 1 -999
box -296 -619 296 619
use sky130_fd_pr__pfet_01v8_lvt_GWB8VV  XM33
timestamp 1739902357
transform 1 0 3684 0 1 -998
box -396 -619 396 619
use sky130_fd_pr__pfet_01v8_lvt_GWB8VV  XM34
timestamp 1739902357
transform 1 0 616 0 1 -999
box -396 -619 396 619
use sky130_fd_pr__nfet_01v8_lvt_VWWV9N  XM35
timestamp 1739902357
transform 1 0 387 0 1 -2360
box -625 -610 625 610
use sky130_fd_pr__nfet_01v8_lvt_VWWV9N  XM36
timestamp 1739902357
transform 1 0 3913 0 1 -2361
box -625 -610 625 610
use sky130_fd_pr__pfet_01v8_lvt_TZF6Y6  XM37
timestamp 1739902357
transform 1 0 4784 0 1 -1245
box -246 -269 246 269
use sky130_fd_pr__nfet_01v8_lvt_PVEEJN  XM38
timestamp 1739902357
transform 1 0 4784 0 1 -2141
box -246 -390 246 390
<< labels >>
flabel metal2 2480 -2065 2680 -1865 0 FreeSans 256 0 0 0 Vin
port 2 nsew
flabel metal1 -254 -3239 -54 -3039 0 FreeSans 256 0 0 0 VGND
port 4 nsew
flabel metal1 162 -348 362 -148 0 FreeSans 256 0 0 0 VPWR
port 0 nsew
flabel metal2 1477 -2065 1677 -1865 0 FreeSans 256 0 0 0 Vref
port 1 nsew
flabel metal2 4884 -1731 5084 -1531 0 FreeSans 256 0 0 0 Vcomp_n
port 3 nsew
<< end >>
