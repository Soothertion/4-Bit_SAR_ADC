magic
tech sky130A
magscale 1 2
timestamp 1739974041
<< nwell >>
rect -625 -619 625 619
<< pmoslvt >>
rect -429 -400 -29 400
rect 29 -400 429 400
<< pdiff >>
rect -487 388 -429 400
rect -487 -388 -475 388
rect -441 -388 -429 388
rect -487 -400 -429 -388
rect -29 388 29 400
rect -29 -388 -17 388
rect 17 -388 29 388
rect -29 -400 29 -388
rect 429 388 487 400
rect 429 -388 441 388
rect 475 -388 487 388
rect 429 -400 487 -388
<< pdiffc >>
rect -475 -388 -441 388
rect -17 -388 17 388
rect 441 -388 475 388
<< nsubdiff >>
rect -589 549 -493 583
rect 493 549 589 583
rect -589 487 -555 549
rect 555 487 589 549
rect -589 -549 -555 -487
rect 555 -549 589 -487
rect -589 -583 -493 -549
rect 493 -583 589 -549
<< nsubdiffcont >>
rect -493 549 493 583
rect -589 -487 -555 487
rect 555 -487 589 487
rect -493 -583 493 -549
<< poly >>
rect -429 481 -29 497
rect -429 447 -413 481
rect -45 447 -29 481
rect -429 400 -29 447
rect 29 481 429 497
rect 29 447 45 481
rect 413 447 429 481
rect 29 400 429 447
rect -429 -447 -29 -400
rect -429 -481 -413 -447
rect -45 -481 -29 -447
rect -429 -497 -29 -481
rect 29 -447 429 -400
rect 29 -481 45 -447
rect 413 -481 429 -447
rect 29 -497 429 -481
<< polycont >>
rect -413 447 -45 481
rect 45 447 413 481
rect -413 -481 -45 -447
rect 45 -481 413 -447
<< locali >>
rect -589 549 -493 583
rect 493 549 589 583
rect -589 487 -555 549
rect 555 487 589 549
rect -429 447 -413 481
rect -45 447 -29 481
rect 29 447 45 481
rect 413 447 429 481
rect -475 388 -441 404
rect -475 -404 -441 -388
rect -17 388 17 404
rect -17 -404 17 -388
rect 441 388 475 404
rect 441 -404 475 -388
rect -429 -481 -413 -447
rect -45 -481 -29 -447
rect 29 -481 45 -447
rect 413 -481 429 -447
rect -589 -549 -555 -487
rect 555 -549 589 -487
rect -589 -583 -493 -549
rect 493 -583 589 -549
<< viali >>
rect -413 447 -45 481
rect 45 447 413 481
rect -475 -388 -441 388
rect -17 -388 17 388
rect 441 -388 475 388
rect -413 -481 -45 -447
rect 45 -481 413 -447
<< metal1 >>
rect -425 481 -33 487
rect -425 447 -413 481
rect -45 447 -33 481
rect -425 441 -33 447
rect 33 481 425 487
rect 33 447 45 481
rect 413 447 425 481
rect 33 441 425 447
rect -481 388 -435 400
rect -481 -388 -475 388
rect -441 -388 -435 388
rect -481 -400 -435 -388
rect -23 388 23 400
rect -23 -388 -17 388
rect 17 -388 23 388
rect -23 -400 23 -388
rect 435 388 481 400
rect 435 -388 441 388
rect 475 -388 481 388
rect 435 -400 481 -388
rect -425 -447 -33 -441
rect -425 -481 -413 -447
rect -45 -481 -33 -447
rect -425 -487 -33 -481
rect 33 -447 425 -441
rect 33 -481 45 -447
rect 413 -481 425 -447
rect 33 -487 425 -481
<< properties >>
string FIXED_BBOX -572 -566 572 566
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 4 l 2.0 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
