magic
tech sky130A
magscale 1 2
timestamp 1739436521
<< pwell >>
rect -246 -271 246 271
<< nmoslvt >>
rect -50 -61 50 61
<< ndiff >>
rect -108 49 -50 61
rect -108 -49 -96 49
rect -62 -49 -50 49
rect -108 -61 -50 -49
rect 50 49 108 61
rect 50 -49 62 49
rect 96 -49 108 49
rect 50 -61 108 -49
<< ndiffc >>
rect -96 -49 -62 49
rect 62 -49 96 49
<< psubdiff >>
rect -210 201 -114 235
rect 114 201 210 235
rect -210 139 -176 201
rect 176 139 210 201
rect -210 -201 -176 -139
rect 176 -201 210 -139
rect -210 -235 -114 -201
rect 114 -235 210 -201
<< psubdiffcont >>
rect -114 201 114 235
rect -210 -139 -176 139
rect 176 -139 210 139
rect -114 -235 114 -201
<< poly >>
rect -50 133 50 149
rect -50 99 -34 133
rect 34 99 50 133
rect -50 61 50 99
rect -50 -99 50 -61
rect -50 -133 -34 -99
rect 34 -133 50 -99
rect -50 -149 50 -133
<< polycont >>
rect -34 99 34 133
rect -34 -133 34 -99
<< locali >>
rect -210 201 -114 235
rect 114 201 210 235
rect -210 139 -176 201
rect 176 139 210 201
rect -50 99 -34 133
rect 34 99 50 133
rect -96 49 -62 65
rect -96 -65 -62 -49
rect 62 49 96 65
rect 62 -65 96 -49
rect -50 -133 -34 -99
rect 34 -133 50 -99
rect -210 -201 -176 -139
rect 176 -201 210 -139
rect -210 -235 -114 -201
rect 114 -235 210 -201
<< viali >>
rect -34 99 34 133
rect -96 -49 -62 49
rect 62 -49 96 49
rect -34 -133 34 -99
<< metal1 >>
rect -46 133 46 139
rect -46 99 -34 133
rect 34 99 46 133
rect -46 93 46 99
rect -102 49 -56 61
rect -102 -49 -96 49
rect -62 -49 -56 49
rect -102 -61 -56 -49
rect 56 49 102 61
rect 56 -49 62 49
rect 96 -49 102 49
rect 56 -61 102 -49
rect -46 -99 46 -93
rect -46 -133 -34 -99
rect 34 -133 46 -99
rect -46 -139 46 -133
<< properties >>
string FIXED_BBOX -193 -218 193 218
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 0.61 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
