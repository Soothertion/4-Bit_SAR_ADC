magic
tech sky130A
magscale 1 2
timestamp 1739902357
<< pwell >>
rect -625 -610 625 610
<< nmoslvt >>
rect -429 -400 -29 400
rect 29 -400 429 400
<< ndiff >>
rect -487 388 -429 400
rect -487 -388 -475 388
rect -441 -388 -429 388
rect -487 -400 -429 -388
rect -29 388 29 400
rect -29 -388 -17 388
rect 17 -388 29 388
rect -29 -400 29 -388
rect 429 388 487 400
rect 429 -388 441 388
rect 475 -388 487 388
rect 429 -400 487 -388
<< ndiffc >>
rect -475 -388 -441 388
rect -17 -388 17 388
rect 441 -388 475 388
<< psubdiff >>
rect -589 540 -493 574
rect 493 540 589 574
rect -589 478 -555 540
rect 555 478 589 540
rect -589 -540 -555 -478
rect 555 -540 589 -478
rect -589 -574 -493 -540
rect 493 -574 589 -540
<< psubdiffcont >>
rect -493 540 493 574
rect -589 -478 -555 478
rect 555 -478 589 478
rect -493 -574 493 -540
<< poly >>
rect -429 472 -29 488
rect -429 438 -413 472
rect -45 438 -29 472
rect -429 400 -29 438
rect 29 472 429 488
rect 29 438 45 472
rect 413 438 429 472
rect 29 400 429 438
rect -429 -438 -29 -400
rect -429 -472 -413 -438
rect -45 -472 -29 -438
rect -429 -488 -29 -472
rect 29 -438 429 -400
rect 29 -472 45 -438
rect 413 -472 429 -438
rect 29 -488 429 -472
<< polycont >>
rect -413 438 -45 472
rect 45 438 413 472
rect -413 -472 -45 -438
rect 45 -472 413 -438
<< locali >>
rect -589 540 -493 574
rect 493 540 589 574
rect -589 478 -555 540
rect 555 478 589 540
rect -429 438 -413 472
rect -45 438 -29 472
rect 29 438 45 472
rect 413 438 429 472
rect -475 388 -441 404
rect -475 -404 -441 -388
rect -17 388 17 404
rect -17 -404 17 -388
rect 441 388 475 404
rect 441 -404 475 -388
rect -429 -472 -413 -438
rect -45 -472 -29 -438
rect 29 -472 45 -438
rect 413 -472 429 -438
rect -589 -540 -555 -478
rect 555 -540 589 -478
rect -589 -574 -493 -540
rect 493 -574 589 -540
<< viali >>
rect -413 438 -45 472
rect 45 438 413 472
rect -475 -388 -441 388
rect -17 -388 17 388
rect 441 -388 475 388
rect -413 -472 -45 -438
rect 45 -472 413 -438
<< metal1 >>
rect -425 472 -33 478
rect -425 438 -413 472
rect -45 438 -33 472
rect -425 432 -33 438
rect 33 472 425 478
rect 33 438 45 472
rect 413 438 425 472
rect 33 432 425 438
rect -481 388 -435 400
rect -481 -388 -475 388
rect -441 -388 -435 388
rect -481 -400 -435 -388
rect -23 388 23 400
rect -23 -388 -17 388
rect 17 -388 23 388
rect -23 -400 23 -388
rect 435 388 481 400
rect 435 -388 441 388
rect 475 -388 481 388
rect 435 -400 481 -388
rect -425 -438 -33 -432
rect -425 -472 -413 -438
rect -45 -472 -33 -438
rect -425 -478 -33 -472
rect 33 -438 425 -432
rect 33 -472 45 -438
rect 413 -472 425 -438
rect 33 -478 425 -472
<< properties >>
string FIXED_BBOX -572 -557 572 557
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 4.0 l 2.0 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
